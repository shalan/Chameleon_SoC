* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[16] IRQ[17] IRQ[18] IRQ[19] IRQ[20] IRQ[21] IRQ[22]
+ IRQ[23] IRQ[24] IRQ[25] IRQ[26] IRQ[27] IRQ[28] IRQ[29] IRQ[30] IRQ[31] MSI_S2 MSI_S3
+ MSO_S2 MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6
+ pwm_S7 scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 VPWR VGND
XFILLER_140_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18869_ _16482_/Y _24157_/Q _16497_/Y _24151_/Q VGND VGND VPWR VPWR _18869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20900_ _20836_/A VGND VGND VPWR VPWR _20900_/X sky130_fd_sc_hd__buf_2
X_21880_ _21880_/A _21867_/Y _21872_/X _21879_/X VGND VGND VPWR VPWR _21880_/X sky130_fd_sc_hd__or4_4
X_20831_ _20831_/A _20831_/B VGND VGND VPWR VPWR _20881_/A sky130_fd_sc_hd__or2_4
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21832__A _22274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22342__A2 _22327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20762_ _13143_/C VGND VGND VPWR VPWR _20768_/B sky130_fd_sc_hd__buf_2
X_23550_ _23582_/CLK _20011_/X VGND VGND VPWR VPWR _20009_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17217__A2_N _17391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16557__B1 _16294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22501_ _22204_/A VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__buf_2
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23481_ _23488_/CLK _23481_/D VGND VGND VPWR VPWR _23481_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20693_ _20693_/A _20693_/B VGND VGND VPWR VPWR _20694_/A sky130_fd_sc_hd__or2_4
XFILLER_167_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22432_ _20864_/Y _22296_/X _20725_/A _21322_/X VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__a2bb2o_4
X_25220_ _25215_/CLK _14170_/X HRESETn VGND VGND VPWR VPWR _14108_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_195_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22363_ _22359_/X _22362_/X _21697_/X VGND VGND VPWR VPWR _22363_/Y sky130_fd_sc_hd__o21ai_4
X_25151_ _24095_/CLK _14413_/X HRESETn VGND VGND VPWR VPWR _20614_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21853__A1 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21314_ _21314_/A VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__buf_2
X_24102_ _25177_/CLK _13655_/Y HRESETn VGND VGND VPWR VPWR _14310_/A sky130_fd_sc_hd__dfrtp_4
X_25082_ _25082_/CLK _14653_/X HRESETn VGND VGND VPWR VPWR _14794_/A sky130_fd_sc_hd__dfrtp_4
X_22294_ _22294_/A _22294_/B VGND VGND VPWR VPWR _22311_/C sky130_fd_sc_hd__nor2_4
X_24033_ _24495_/CLK _20778_/X HRESETn VGND VGND VPWR VPWR _24033_/Q sky130_fd_sc_hd__dfrtp_4
X_21245_ _14687_/A VGND VGND VPWR VPWR _21246_/A sky130_fd_sc_hd__inv_2
XANTENNA__25098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21176_ _16454_/Y _21574_/A _16379_/A _21175_/X VGND VGND VPWR VPWR _21177_/C sky130_fd_sc_hd__a211o_4
XFILLER_89_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20127_ _19859_/X _13757_/X VGND VGND VPWR VPWR _20128_/A sky130_fd_sc_hd__and2_4
XFILLER_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20058_ _13762_/X _14706_/A _13774_/X _13775_/X VGND VGND VPWR VPWR _20059_/A sky130_fd_sc_hd__or4_4
X_24935_ _24354_/CLK _15543_/X HRESETn VGND VGND VPWR VPWR _11731_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11900_ _11900_/A VGND VGND VPWR VPWR _11901_/A sky130_fd_sc_hd__inv_2
XANTENNA__19982__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12880_ _12790_/A _12880_/B VGND VGND VPWR VPWR _12880_/X sky130_fd_sc_hd__or2_4
X_24866_ _24867_/CLK _24866_/D HRESETn VGND VGND VPWR VPWR _24866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_128_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _24258_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11830_/X VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__buf_2
X_23817_ _23454_/CLK _23817_/D VGND VGND VPWR VPWR _13312_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24799_/CLK _15910_/X HRESETn VGND VGND VPWR VPWR _22428_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22557__B _16382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14550_ _14550_/A _14550_/B VGND VGND VPWR VPWR _14550_/X sky130_fd_sc_hd__or2_4
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24662__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _25553_/Q VGND VGND VPWR VPWR _11762_/Y sky130_fd_sc_hd__inv_2
X_23748_ _23669_/CLK _23748_/D VGND VGND VPWR VPWR _17963_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13500_/Y _13498_/X _11871_/X _13498_/X VGND VGND VPWR VPWR _13501_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _25127_/Q VGND VGND VPWR VPWR _14481_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11691_/A _24232_/Q _13690_/A _11692_/Y VGND VGND VPWR VPWR _11693_/X sky130_fd_sc_hd__o22a_4
X_23679_ _23582_/CLK _23679_/D VGND VGND VPWR VPWR _19641_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16219_/Y _16215_/X _15960_/X _16215_/X VGND VGND VPWR VPWR _16220_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13243_/X _13432_/B VGND VGND VPWR VPWR _13432_/X sky130_fd_sc_hd__or2_4
X_25418_ _25410_/CLK _12709_/Y HRESETn VGND VGND VPWR VPWR _12574_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _16150_/Y _16148_/X _15905_/X _16148_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__a2bb2o_4
X_13363_ _13242_/X _13361_/X _13363_/C VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__and3_4
X_25349_ _25368_/CLK _13102_/X HRESETn VGND VGND VPWR VPWR _25349_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16571__A _16571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15102_ _15396_/A _24585_/Q _15396_/A _24585_/Q VGND VGND VPWR VPWR _15102_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12314_ _24835_/Q VGND VGND VPWR VPWR _12314_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16082_ _24722_/Q VGND VGND VPWR VPWR _16082_/Y sky130_fd_sc_hd__inv_2
X_13294_ _13241_/X _13289_/X _13293_/X VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__or3_4
XFILLER_154_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15033_ _15282_/A _15000_/Y _25023_/Q _15032_/Y VGND VGND VPWR VPWR _15033_/X sky130_fd_sc_hd__a2bb2o_4
X_19910_ _19904_/Y VGND VGND VPWR VPWR _19910_/X sky130_fd_sc_hd__buf_2
XFILLER_6_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12245_ _12439_/B _22644_/A _12296_/B _22644_/A VGND VGND VPWR VPWR _12245_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12176_ _25475_/Q _14334_/A _12175_/X _12170_/X VGND VGND VPWR VPWR _12177_/A sky130_fd_sc_hd__a211o_4
X_19841_ _23611_/Q VGND VGND VPWR VPWR _22230_/B sky130_fd_sc_hd__inv_2
X_16984_ _24729_/Q _24386_/Q _16063_/Y _17142_/A VGND VGND VPWR VPWR _16984_/X sky130_fd_sc_hd__o22a_4
X_19772_ HWDATA[5] VGND VGND VPWR VPWR _19772_/X sky130_fd_sc_hd__buf_2
XFILLER_122_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15935_ _15664_/X _15844_/X _15933_/X _24786_/Q _15934_/X VGND VGND VPWR VPWR _24786_/D
+ sky130_fd_sc_hd__a32o_4
X_18723_ _18722_/X VGND VGND VPWR VPWR _18723_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11848__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_24_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22572__A2 _22571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18654_ _24154_/Q VGND VGND VPWR VPWR _18744_/A sky130_fd_sc_hd__buf_2
X_15866_ _21173_/B VGND VGND VPWR VPWR _15866_/X sky130_fd_sc_hd__buf_2
XFILLER_237_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_87_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14817_ _14817_/A VGND VGND VPWR VPWR _14835_/A sky130_fd_sc_hd__buf_2
X_17605_ _17604_/X VGND VGND VPWR VPWR _17606_/B sky130_fd_sc_hd__inv_2
X_18585_ _18493_/A VGND VGND VPWR VPWR _18598_/C sky130_fd_sc_hd__buf_2
XFILLER_224_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15797_ _15796_/X VGND VGND VPWR VPWR _15797_/X sky130_fd_sc_hd__buf_2
XFILLER_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20828__A1_N _20698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17536_ _25542_/Q _17578_/B _11849_/Y _17538_/A VGND VGND VPWR VPWR _17542_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15650__A _22121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14748_ _14740_/X _14747_/Y _14734_/A _14732_/Y VGND VGND VPWR VPWR _14748_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ _17465_/X VGND VGND VPWR VPWR _17467_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14679_ _13628_/B _14679_/B VGND VGND VPWR VPWR _19436_/B sky130_fd_sc_hd__or2_4
XFILLER_177_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16418_ _15127_/Y _16415_/X _16417_/X _16415_/X VGND VGND VPWR VPWR _16418_/X sky130_fd_sc_hd__a2bb2o_4
X_19206_ _19205_/Y _19203_/X _19184_/X _19203_/X VGND VGND VPWR VPWR _23830_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17398_ _17398_/A _17398_/B VGND VGND VPWR VPWR _17399_/B sky130_fd_sc_hd__or2_4
XANTENNA__22483__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19137_ _19136_/Y _19134_/X _19048_/X _19134_/X VGND VGND VPWR VPWR _19137_/X sky130_fd_sc_hd__a2bb2o_4
X_16349_ HWDATA[10] VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__buf_2
XFILLER_145_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19068_ _19061_/A VGND VGND VPWR VPWR _19068_/X sky130_fd_sc_hd__buf_2
XFILLER_218_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21099__A _23087_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18019_ _18060_/A _23851_/Q VGND VGND VPWR VPWR _18022_/B sky130_fd_sc_hd__or2_4
XANTENNA__13525__B1 _13524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12328__B2 _12327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21030_ _22306_/A VGND VGND VPWR VPWR _21060_/A sky130_fd_sc_hd__buf_2
XANTENNA__25191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21827__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20271__B1 _20249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11839__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22981_ _21449_/A VGND VGND VPWR VPWR _23117_/A sky130_fd_sc_hd__buf_2
XFILLER_228_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24720_ _23386_/CLK _24720_/D HRESETn VGND VGND VPWR VPWR _21071_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13345__A _13212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21932_ _18314_/X VGND VGND VPWR VPWR _21938_/A sky130_fd_sc_hd__buf_2
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24651_ _24651_/CLK _24651_/D HRESETn VGND VGND VPWR VPWR _21021_/A sky130_fd_sc_hd__dfrtp_4
X_21863_ _21858_/X _21863_/B _21860_/X _21863_/D VGND VGND VPWR VPWR _21863_/X sky130_fd_sc_hd__and4_4
XANTENNA__19716__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23602_ _25068_/CLK _19868_/X VGND VGND VPWR VPWR _23602_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15560__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20814_ _24042_/Q _20810_/X _20818_/B VGND VGND VPWR VPWR _20814_/Y sky130_fd_sc_hd__a21oi_4
X_21794_ _22237_/A _21794_/B _21793_/X VGND VGND VPWR VPWR _21794_/X sky130_fd_sc_hd__or3_4
X_24582_ _24562_/CLK _24582_/D HRESETn VGND VGND VPWR VPWR _16472_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23582_/CLK _23533_/D VGND VGND VPWR VPWR _23533_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20745_ _20739_/X _20741_/Y _24908_/Q _20744_/X VGND VGND VPWR VPWR _20745_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20676_ _23999_/Q _17408_/B _17410_/A VGND VGND VPWR VPWR _20676_/Y sky130_fd_sc_hd__a21oi_4
X_23464_ _23466_/CLK _23464_/D VGND VGND VPWR VPWR _18114_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23276__B1 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25203_ _25204_/CLK _14241_/X HRESETn VGND VGND VPWR VPWR _25203_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22415_ _25532_/Q _22411_/X _21042_/X _22414_/X VGND VGND VPWR VPWR _22415_/X sky130_fd_sc_hd__a211o_4
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23395_ _23395_/CLK _20421_/X VGND VGND VPWR VPWR _23395_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25134_ _25148_/CLK _25134_/D HRESETn VGND VGND VPWR VPWR _14103_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22346_ _21941_/A _22346_/B VGND VGND VPWR VPWR _22348_/B sky130_fd_sc_hd__or2_4
XANTENNA__16702__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22277_ _22277_/A VGND VGND VPWR VPWR _22277_/Y sky130_fd_sc_hd__inv_2
X_25065_ _24258_/CLK _14784_/X HRESETn VGND VGND VPWR VPWR _25065_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23043__A3 _22291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12030_ _12030_/A VGND VGND VPWR VPWR _12030_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21228_ _15650_/X VGND VGND VPWR VPWR _22808_/A sky130_fd_sc_hd__buf_2
X_24016_ _24015_/CLK _20703_/Y HRESETn VGND VGND VPWR VPWR _13131_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18455__B1 _16271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15728__A1_N _12555_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21159_ _21158_/Y _21353_/A _14890_/Y _14442_/A VGND VGND VPWR VPWR _21164_/B sky130_fd_sc_hd__o22a_4
XFILLER_120_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13981_ scl_oen_o_S5 _13975_/X _13976_/Y _13980_/Y VGND VGND VPWR VPWR _13982_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15720_ _15719_/X VGND VGND VPWR VPWR _15720_/X sky130_fd_sc_hd__buf_2
XANTENNA__22554__A2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ _12931_/X VGND VGND VPWR VPWR _25389_/D sky130_fd_sc_hd__inv_2
X_24918_ _24915_/CLK _24918_/D HRESETn VGND VGND VPWR VPWR _24918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16769__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24843__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15651_ _14386_/A _15650_/X VGND VGND VPWR VPWR _15651_/X sky130_fd_sc_hd__or2_4
XFILLER_218_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12863_ _12765_/Y _12862_/X VGND VGND VPWR VPWR _12863_/X sky130_fd_sc_hd__or2_4
X_24849_ _24849_/CLK _24849_/D HRESETn VGND VGND VPWR VPWR _24849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19707__B1 _19560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14577_/X _14595_/X _14601_/Y _14599_/X _25097_/Q VGND VGND VPWR VPWR _14602_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11803_/X VGND VGND VPWR VPWR _11814_/X sky130_fd_sc_hd__buf_2
X_18370_ _18370_/A _18360_/Y VGND VGND VPWR VPWR _18370_/Y sky130_fd_sc_hd__nor2_4
XFILLER_33_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15581_/Y _15577_/X _11770_/X _15577_/X VGND VGND VPWR VPWR _15582_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15992__A1 _15797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _22490_/A VGND VGND VPWR VPWR _12794_/Y sky130_fd_sc_hd__inv_2
XPHY_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17186_/A _17321_/B VGND VGND VPWR VPWR _17321_/X sky130_fd_sc_hd__or2_4
XPHY_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _25111_/Q _14520_/X _25110_/Q _14522_/X VGND VGND VPWR VPWR _14533_/X sky130_fd_sc_hd__o22a_4
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11744_/X VGND VGND VPWR VPWR _22575_/A sky130_fd_sc_hd__buf_2
XFILLER_159_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17194__B1 _16354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17362_/A _17358_/C _17357_/A _17252_/D VGND VGND VPWR VPWR _17252_/X sky130_fd_sc_hd__or4_4
XFILLER_159_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14464_ _20608_/A _14463_/X _14420_/X _14463_/X VGND VGND VPWR VPWR _25134_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11676_/A VGND VGND VPWR VPWR _11676_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22195__A2_N _22176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _16227_/A VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__buf_2
X_13415_ _13310_/X _13413_/X _13415_/C VGND VGND VPWR VPWR _13415_/X sky130_fd_sc_hd__and3_4
XFILLER_186_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17183_ _17183_/A VGND VGND VPWR VPWR _17184_/A sky130_fd_sc_hd__inv_2
X_14395_ _14395_/A VGND VGND VPWR VPWR _14395_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23282__A3 _22861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16134_ _22792_/A VGND VGND VPWR VPWR _16134_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13346_ _13410_/A _13346_/B VGND VGND VPWR VPWR _13346_/X sky130_fd_sc_hd__or2_4
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16065_ _16065_/A VGND VGND VPWR VPWR _16065_/Y sky130_fd_sc_hd__inv_2
X_13277_ _13315_/A _13277_/B _13276_/X VGND VGND VPWR VPWR _13285_/B sky130_fd_sc_hd__or3_4
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15016_ _15016_/A VGND VGND VPWR VPWR _15268_/A sky130_fd_sc_hd__buf_2
X_12228_ _12228_/A VGND VGND VPWR VPWR _12228_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18446__B1 _23250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19824_ _23617_/Q VGND VGND VPWR VPWR _19824_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12159_ _12113_/Y _12158_/X _12113_/Y _12158_/X VGND VGND VPWR VPWR _12166_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19755_ _13401_/B VGND VGND VPWR VPWR _19755_/Y sky130_fd_sc_hd__inv_2
X_16967_ _16055_/Y _24389_/Q _16055_/Y _24389_/Q VGND VGND VPWR VPWR _16967_/X sky130_fd_sc_hd__a2bb2o_4
X_18706_ _18705_/X VGND VGND VPWR VPWR _18708_/B sky130_fd_sc_hd__inv_2
XFILLER_209_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17860__A _16920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15918_ _15714_/X _15902_/X _15851_/X _24790_/Q _15871_/X VGND VGND VPWR VPWR _15918_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24584__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16898_ _16896_/Y _16889_/X _16897_/X _14791_/X VGND VGND VPWR VPWR _16898_/X sky130_fd_sc_hd__a2bb2o_4
X_19686_ _13361_/B VGND VGND VPWR VPWR _19686_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15849_ _12353_/Y _15842_/X _15848_/X _15818_/A VGND VGND VPWR VPWR _15849_/X sky130_fd_sc_hd__a2bb2o_4
X_18637_ _24140_/Q VGND VGND VPWR VPWR _18637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16476__A _16495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_111_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24495_/CLK sky130_fd_sc_hd__clkbuf_1
X_18568_ _18482_/A _18567_/X VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__or2_4
XFILLER_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_174_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _23871_/CLK sky130_fd_sc_hd__clkbuf_1
X_17519_ _25533_/Q _24304_/Q _11837_/Y _17518_/Y VGND VGND VPWR VPWR _17524_/B sky130_fd_sc_hd__o22a_4
X_18499_ _18499_/A VGND VGND VPWR VPWR _18500_/B sky130_fd_sc_hd__inv_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20530_ _20530_/A _20456_/X VGND VGND VPWR VPWR _20531_/D sky130_fd_sc_hd__and2_4
XFILLER_220_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19813__A2_N _19806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15735__A1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20461_ _20444_/A _20609_/B _20461_/C _20461_/D VGND VGND VPWR VPWR _20461_/X sky130_fd_sc_hd__and4_4
X_22200_ _21235_/X VGND VGND VPWR VPWR _22425_/B sky130_fd_sc_hd__buf_2
XANTENNA__25372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23180_ _23136_/X _23180_/B VGND VGND VPWR VPWR _23180_/Y sky130_fd_sc_hd__nor2_4
XFILLER_229_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20392_ _22045_/B _20386_/X _19632_/A _20391_/X VGND VGND VPWR VPWR _23409_/D sky130_fd_sc_hd__a2bb2o_4
X_22131_ _22131_/A VGND VGND VPWR VPWR _22131_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22769__C1 _22768_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22062_ _22062_/A _23354_/B VGND VGND VPWR VPWR _22062_/Y sky130_fd_sc_hd__nand2_4
XFILLER_160_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21013_ _21012_/Y _23983_/Q _21013_/C VGND VGND VPWR VPWR _23981_/D sky130_fd_sc_hd__and3_4
XANTENNA__20244__B1 _20243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15555__A _16003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22964_ _16679_/Y _22808_/A _15596_/Y _22845_/X VGND VGND VPWR VPWR _22964_/X sky130_fd_sc_hd__o22a_4
XFILLER_244_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18204__A3 _18203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22388__A _22388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24703_ _25444_/CLK _16133_/X HRESETn VGND VGND VPWR VPWR _24703_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21915_ _14766_/X _19933_/Y VGND VGND VPWR VPWR _21915_/X sky130_fd_sc_hd__or2_4
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_70_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22895_ _23008_/A _22894_/X VGND VGND VPWR VPWR _22895_/Y sky130_fd_sc_hd__nor2_4
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14226__B2 _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24634_ _24629_/CLK _16330_/X HRESETn VGND VGND VPWR VPWR _24634_/Q sky130_fd_sc_hd__dfrtp_4
X_21846_ _13135_/A _21844_/X _24902_/Q _22695_/B VGND VGND VPWR VPWR _21846_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24565_ _24542_/CLK _16516_/X HRESETn VGND VGND VPWR VPWR _24565_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ _14709_/X _21769_/X _21776_/X VGND VGND VPWR VPWR _21777_/X sky130_fd_sc_hd__or3_4
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23516_ _23516_/CLK _20103_/X VGND VGND VPWR VPWR _20099_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_196_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20728_ _15628_/Y _20716_/X _20724_/X _20727_/Y VGND VGND VPWR VPWR _20728_/X sky130_fd_sc_hd__o22a_4
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24496_ _24532_/CLK _16700_/X HRESETn VGND VGND VPWR VPWR _16699_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_184_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20636__A _14816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23447_ _24295_/CLK _20292_/X VGND VGND VPWR VPWR _23447_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20659_ _20659_/A VGND VGND VPWR VPWR _20659_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ _13200_/A _13198_/X _13199_/X VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__and3_4
X_14180_ _14190_/A _23968_/Q VGND VGND VPWR VPWR _14181_/A sky130_fd_sc_hd__or2_4
X_23378_ _23378_/A VGND VGND VPWR VPWR IRQ[22] sky130_fd_sc_hd__buf_2
XANTENNA__25042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13131_ _13131_/A _13131_/B VGND VGND VPWR VPWR _13132_/B sky130_fd_sc_hd__nor2_4
X_25117_ _24095_/CLK _14513_/X HRESETn VGND VGND VPWR VPWR _25117_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22329_ _21040_/Y _22328_/X VGND VGND VPWR VPWR _22329_/X sky130_fd_sc_hd__and2_4
XFILLER_180_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13062_ _12997_/C _13074_/A VGND VGND VPWR VPWR _13066_/B sky130_fd_sc_hd__or2_4
X_25048_ _24000_/CLK _25048_/D HRESETn VGND VGND VPWR VPWR _14873_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12013_ _12001_/X VGND VGND VPWR VPWR _12013_/Y sky130_fd_sc_hd__inv_2
X_17870_ _17872_/B VGND VGND VPWR VPWR _17871_/B sky130_fd_sc_hd__inv_2
XANTENNA__21983__B1 _13793_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16821_ _14928_/Y _16816_/X HWDATA[24] _16820_/X VGND VGND VPWR VPWR _16821_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16752_ _16762_/A VGND VGND VPWR VPWR _16752_/X sky130_fd_sc_hd__buf_2
X_19540_ _23711_/Q VGND VGND VPWR VPWR _21692_/B sky130_fd_sc_hd__inv_2
XFILLER_171_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13964_ _13964_/A _13948_/C _15435_/B VGND VGND VPWR VPWR _13969_/A sky130_fd_sc_hd__or3_4
XANTENNA__21735__B1 _15482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22298__A _22298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15703_ _15703_/A VGND VGND VPWR VPWR _15703_/X sky130_fd_sc_hd__buf_2
XFILLER_207_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12915_ _12917_/B VGND VGND VPWR VPWR _12915_/Y sky130_fd_sc_hd__inv_2
X_16683_ _16682_/Y _16680_/X _16414_/X _16680_/X VGND VGND VPWR VPWR _24503_/D sky130_fd_sc_hd__a2bb2o_4
X_19471_ _19470_/Y _19466_/X _19402_/X _19466_/X VGND VGND VPWR VPWR _19471_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25136__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13895_ _24005_/Q VGND VGND VPWR VPWR _13976_/A sky130_fd_sc_hd__buf_2
XFILLER_47_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15634_ _15634_/A VGND VGND VPWR VPWR _15634_/Y sky130_fd_sc_hd__inv_2
X_18422_ _16201_/A _24192_/Q _16201_/Y _18488_/B VGND VGND VPWR VPWR _18429_/A sky130_fd_sc_hd__o22a_4
XANTENNA__25199__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12846_ _12846_/A _12845_/X VGND VGND VPWR VPWR _12846_/X sky130_fd_sc_hd__or2_4
XFILLER_221_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12779__A1 _25381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18353_ _13200_/A _18351_/X _18352_/Y VGND VGND VPWR VPWR _18353_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12779__B2 _12778_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21930__A _21212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15565_ _21855_/B VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_247_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24975_/CLK sky130_fd_sc_hd__clkbuf_1
X_12777_ _12777_/A VGND VGND VPWR VPWR _12777_/X sky130_fd_sc_hd__buf_2
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22160__B1 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17304_ _24371_/Q _17303_/Y VGND VGND VPWR VPWR _17304_/X sky130_fd_sc_hd__or2_4
XFILLER_203_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14514_/X _14515_/Y _14510_/B VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__a21o_4
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _14385_/A _16190_/B _16378_/C _15791_/D VGND VGND VPWR VPWR _11728_/X sky130_fd_sc_hd__or4_4
X_18284_ _17733_/A VGND VGND VPWR VPWR _18285_/D sky130_fd_sc_hd__buf_2
XFILLER_30_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15496_ _20437_/A _15495_/X VGND VGND VPWR VPWR _15496_/X sky130_fd_sc_hd__or2_4
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17235_ _16293_/Y _17244_/A _16293_/Y _17244_/A VGND VGND VPWR VPWR _17235_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _14441_/Y _14446_/X _14420_/X _14446_/X VGND VGND VPWR VPWR _14447_/X sky130_fd_sc_hd__a2bb2o_4
X_11659_ _11712_/A VGND VGND VPWR VPWR _11660_/A sky130_fd_sc_hd__inv_2
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17166_ _17048_/Y _17166_/B VGND VGND VPWR VPWR _17167_/B sky130_fd_sc_hd__or2_4
XFILLER_128_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14378_ _14364_/A _14377_/X _12094_/A _14369_/X VGND VGND VPWR VPWR _14378_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22463__B2 _16552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16117_ _16115_/Y _16111_/X _15957_/X _16116_/X VGND VGND VPWR VPWR _24710_/D sky130_fd_sc_hd__a2bb2o_4
X_13329_ _13468_/A _13329_/B VGND VGND VPWR VPWR _13329_/X sky130_fd_sc_hd__or2_4
XFILLER_171_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17097_ _17393_/B _17094_/B _17097_/C VGND VGND VPWR VPWR _17097_/X sky130_fd_sc_hd__or3_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12586__A2_N _24875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16048_ _24735_/Q VGND VGND VPWR VPWR _16048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21377__A _21369_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21423__C1 _21422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19092__B1 _19091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24765__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17188__A1_N _24638_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19807_ _16887_/X VGND VGND VPWR VPWR _19807_/X sky130_fd_sc_hd__buf_2
XFILLER_85_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17999_ _18189_/A _19463_/A VGND VGND VPWR VPWR _18002_/B sky130_fd_sc_hd__or2_4
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19738_ _13464_/B VGND VGND VPWR VPWR _19738_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19669_ _13429_/B VGND VGND VPWR VPWR _19669_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15405__B1 _15348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21700_ _21679_/X _21699_/X _21511_/X VGND VGND VPWR VPWR _21700_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22680_ _22680_/A _22678_/X _22679_/X _22294_/A VGND VGND VPWR VPWR _22681_/A sky130_fd_sc_hd__and4_4
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19122__A2_N _19121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21631_ _21627_/X _21630_/X _14758_/X VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24350_ _24354_/CLK _24350_/D HRESETn VGND VGND VPWR VPWR _17250_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12539__A2_N _24860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25553__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21562_ _14402_/Y _14203_/X _14474_/Y _17424_/X VGND VGND VPWR VPWR _21563_/D sky130_fd_sc_hd__o22a_4
X_23301_ _17270_/C _22493_/X _25403_/Q _22453_/X VGND VGND VPWR VPWR _23301_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20513_ _14073_/A _20457_/X VGND VGND VPWR VPWR _20513_/X sky130_fd_sc_hd__and2_4
XFILLER_138_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21493_ _21493_/A _21490_/X _21493_/C VGND VGND VPWR VPWR _21493_/X sky130_fd_sc_hd__and3_4
X_24281_ _24283_/CLK _24281_/D HRESETn VGND VGND VPWR VPWR _24281_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20444_ _20444_/A _24098_/Q VGND VGND VPWR VPWR _20446_/C sky130_fd_sc_hd__or2_4
X_23232_ _23052_/X _23231_/X _22484_/X _12591_/A _23120_/X VGND VGND VPWR VPWR _23233_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18658__B1 _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20375_ _20374_/Y _20370_/X _19639_/A _20370_/X VGND VGND VPWR VPWR _20375_/X sky130_fd_sc_hd__a2bb2o_4
X_23163_ _23052_/X _23162_/X _22986_/X _24886_/Q _23120_/X VGND VGND VPWR VPWR _23164_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22114_ _22113_/X VGND VGND VPWR VPWR _22114_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23094_ _12780_/Y _21890_/X _17753_/B _22839_/X VGND VGND VPWR VPWR _23094_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15892__B1 _11797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22045_ _22034_/A _22045_/B VGND VGND VPWR VPWR _22045_/X sky130_fd_sc_hd__or2_4
XANTENNA__19083__B1 _19012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15644__B1 _15486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23996_ _23998_/CLK _20667_/Y HRESETn VGND VGND VPWR VPWR _17405_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22947_ _22947_/A VGND VGND VPWR VPWR _22947_/X sky130_fd_sc_hd__buf_2
XFILLER_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12700_ _12700_/A VGND VGND VPWR VPWR _12700_/Y sky130_fd_sc_hd__inv_2
X_13680_ _13680_/A VGND VGND VPWR VPWR _13680_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22878_ _24635_/Q _22789_/B VGND VGND VPWR VPWR _22878_/X sky130_fd_sc_hd__or2_4
XFILLER_232_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12631_ _12642_/A _12642_/B _12631_/C _12642_/D VGND VGND VPWR VPWR _12631_/X sky130_fd_sc_hd__or4_4
X_24617_ _24485_/CLK _24617_/D HRESETn VGND VGND VPWR VPWR _24617_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21829_ _21468_/X _19638_/Y VGND VGND VPWR VPWR _21830_/C sky130_fd_sc_hd__or2_4
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _15303_/A _15352_/B _15349_/Y VGND VGND VPWR VPWR _25006_/D sky130_fd_sc_hd__o21a_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19220__A _19085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_0_0_HCLK clkbuf_7_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_12562_ _25408_/Q _12561_/A _12742_/A _12561_/Y VGND VGND VPWR VPWR _12566_/C sky130_fd_sc_hd__o22a_4
X_24548_ _24542_/CLK _16563_/X HRESETn VGND VGND VPWR VPWR _16562_/A sky130_fd_sc_hd__dfrtp_4
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15591__A1_N _15588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_14_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23799_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _14300_/X VGND VGND VPWR VPWR _14301_/Y sky130_fd_sc_hd__inv_2
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _15281_/A VGND VGND VPWR VPWR _15282_/B sky130_fd_sc_hd__inv_2
XFILLER_12_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12501_/A _12491_/X _12493_/C VGND VGND VPWR VPWR _25447_/D sky130_fd_sc_hd__and3_4
X_24479_ _24473_/CLK _24479_/D HRESETn VGND VGND VPWR VPWR _24479_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_77_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24781_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17020_ _17020_/A _17015_/X _17020_/C _17020_/D VGND VGND VPWR VPWR _17026_/C sky130_fd_sc_hd__or4_4
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _14232_/A _14232_/B VGND VGND VPWR VPWR _14233_/A sky130_fd_sc_hd__nor2_4
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22445__A1 _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18649__B1 _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14163_ _14162_/X VGND VGND VPWR VPWR _14163_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13114_ _13114_/A VGND VGND VPWR VPWR _13114_/Y sky130_fd_sc_hd__inv_2
X_14094_ _14028_/A _14090_/X _14087_/X _14027_/B _14093_/X VGND VGND VPWR VPWR _25237_/D
+ sky130_fd_sc_hd__a32o_4
X_18971_ _13354_/B VGND VGND VPWR VPWR _18971_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22748__A2 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _13038_/B VGND VGND VPWR VPWR _13046_/B sky130_fd_sc_hd__inv_2
X_17922_ _13551_/X _14778_/X _14628_/Y VGND VGND VPWR VPWR _17922_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12612__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17853_ _17763_/Y _17847_/X _17798_/X _17849_/Y VGND VGND VPWR VPWR _17853_/X sky130_fd_sc_hd__a211o_4
X_16804_ _16552_/A _16382_/B VGND VGND VPWR VPWR _16857_/A sky130_fd_sc_hd__nor2_4
XANTENNA__24105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14996_ _14996_/A VGND VGND VPWR VPWR _14996_/X sky130_fd_sc_hd__buf_2
X_17784_ _17784_/A VGND VGND VPWR VPWR _17784_/Y sky130_fd_sc_hd__inv_2
X_19523_ _21467_/B _19520_/X _11964_/X _19520_/X VGND VGND VPWR VPWR _19523_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13947_ _13958_/A _13942_/X VGND VGND VPWR VPWR _13947_/Y sky130_fd_sc_hd__nand2_4
X_16735_ _15337_/A _16734_/X _16729_/X _16734_/X VGND VGND VPWR VPWR _16735_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13443__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16666_ _16666_/A VGND VGND VPWR VPWR _16666_/Y sky130_fd_sc_hd__inv_2
X_19454_ _19048_/A VGND VGND VPWR VPWR _19454_/X sky130_fd_sc_hd__buf_2
X_13878_ _25255_/Q _13870_/X _22129_/A _13872_/X VGND VGND VPWR VPWR _13878_/X sky130_fd_sc_hd__o22a_4
XFILLER_179_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15617_ _22651_/A _15614_/X _11822_/X _15614_/X VGND VGND VPWR VPWR _15617_/X sky130_fd_sc_hd__a2bb2o_4
X_18405_ _24173_/Q VGND VGND VPWR VPWR _18479_/D sky130_fd_sc_hd__inv_2
XFILLER_201_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12829_ _23231_/A VGND VGND VPWR VPWR _12829_/Y sky130_fd_sc_hd__inv_2
X_16597_ _16618_/A VGND VGND VPWR VPWR _16597_/X sky130_fd_sc_hd__buf_2
X_19385_ _19385_/A VGND VGND VPWR VPWR _19385_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15548_ _17448_/B _15544_/X HADDR[2] _15547_/X VGND VGND VPWR VPWR _15548_/X sky130_fd_sc_hd__a2bb2o_4
X_18336_ _17477_/A _18937_/B _17477_/B VGND VGND VPWR VPWR _19119_/C sky130_fd_sc_hd__or3_4
XFILLER_188_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18267_ _18267_/A VGND VGND VPWR VPWR _23358_/A sky130_fd_sc_hd__inv_2
XANTENNA__21892__C1 _21113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15479_ _15479_/A VGND VGND VPWR VPWR _15479_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17218_ _16343_/Y _17258_/A _16343_/Y _17258_/A VGND VGND VPWR VPWR _17218_/X sky130_fd_sc_hd__a2bb2o_4
X_18198_ _18166_/A _18198_/B _18198_/C VGND VGND VPWR VPWR _18202_/B sky130_fd_sc_hd__and3_4
XFILLER_175_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17149_ _16992_/Y _17142_/X VGND VGND VPWR VPWR _17149_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20160_ _23496_/Q VGND VGND VPWR VPWR _21790_/B sky130_fd_sc_hd__inv_2
XANTENNA__14677__B2 _13610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15874__B1 _23290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20091_ _20090_/Y _20086_/X _19753_/X _20086_/X VGND VGND VPWR VPWR _20091_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17508__A2_N _24312_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15833__A _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23850_ _23850_/CLK _19153_/X VGND VGND VPWR VPWR _19150_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19305__A _19148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22801_ _22476_/A VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__buf_2
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23781_ _24252_/CLK _23781_/D VGND VGND VPWR VPWR _18209_/B sky130_fd_sc_hd__dfxtp_4
X_20993_ _24129_/Q _24127_/Q _24128_/Q _20992_/X VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__o22a_4
XFILLER_225_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25520_ _25520_/CLK _25520_/D HRESETn VGND VGND VPWR VPWR _17711_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__12895__C _12609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22732_ _22732_/A VGND VGND VPWR VPWR _23106_/A sky130_fd_sc_hd__buf_2
XFILLER_169_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18439__A1_N _16244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25451_ _25454_/CLK _25451_/D HRESETn VGND VGND VPWR VPWR _12250_/A sky130_fd_sc_hd__dfrtp_4
X_22663_ _15718_/A _22662_/X _22148_/C _16051_/A _16003_/A VGND VGND VPWR VPWR _22663_/X
+ sky130_fd_sc_hd__a32o_4
X_24402_ _24952_/CLK _17092_/X HRESETn VGND VGND VPWR VPWR _24402_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21614_ _21644_/A _19850_/Y VGND VGND VPWR VPWR _21617_/B sky130_fd_sc_hd__or2_4
XFILLER_240_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25382_ _25402_/CLK _12965_/X HRESETn VGND VGND VPWR VPWR _12793_/A sky130_fd_sc_hd__dfrtp_4
X_22594_ _13553_/Y _22706_/B VGND VGND VPWR VPWR _22594_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_230_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _25200_/CLK sky130_fd_sc_hd__clkbuf_1
X_24333_ _24334_/CLK _24333_/D HRESETn VGND VGND VPWR VPWR _17440_/A sky130_fd_sc_hd__dfrtp_4
X_21545_ _15565_/X _21544_/X _21445_/X _24827_/Q _21341_/X VGND VGND VPWR VPWR _21545_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13800__B _14264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24264_ _24715_/CLK _17894_/X HRESETn VGND VGND VPWR VPWR _16935_/A sky130_fd_sc_hd__dfrtp_4
X_21476_ _21476_/A VGND VGND VPWR VPWR _21673_/A sky130_fd_sc_hd__buf_2
XFILLER_181_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23215_ _23136_/X _23215_/B VGND VGND VPWR VPWR _23215_/Y sky130_fd_sc_hd__nor2_4
X_20427_ _13278_/B VGND VGND VPWR VPWR _20427_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24195_ _24651_/CLK _24195_/D HRESETn VGND VGND VPWR VPWR _21109_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24687__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23146_ _23249_/A _23145_/X VGND VGND VPWR VPWR _23146_/Y sky130_fd_sc_hd__nor2_4
X_20358_ _23421_/Q VGND VGND VPWR VPWR _21991_/B sky130_fd_sc_hd__inv_2
XANTENNA__24616__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20289_ _21787_/B _20284_/X _19803_/A _20284_/X VGND VGND VPWR VPWR _23448_/D sky130_fd_sc_hd__a2bb2o_4
X_23077_ _24575_/Q _22897_/X _22816_/X VGND VGND VPWR VPWR _23077_/X sky130_fd_sc_hd__o21a_4
X_22028_ _22028_/A _20043_/Y VGND VGND VPWR VPWR _22029_/C sky130_fd_sc_hd__or2_4
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15617__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14850_ _25056_/Q _14811_/B _25056_/Q _14811_/B VGND VGND VPWR VPWR _14850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13801_ _18268_/A VGND VGND VPWR VPWR _13802_/A sky130_fd_sc_hd__inv_2
X_14781_ _14781_/A _14781_/B _14778_/X _14780_/X VGND VGND VPWR VPWR _14781_/X sky130_fd_sc_hd__or4_4
X_11993_ _11981_/X VGND VGND VPWR VPWR _11993_/Y sky130_fd_sc_hd__inv_2
X_23979_ _24979_/CLK _23979_/D HRESETn VGND VGND VPWR VPWR _23979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22363__B1 _21697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16520_ _16533_/A VGND VGND VPWR VPWR _16520_/X sky130_fd_sc_hd__buf_2
XFILLER_205_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13732_ _11685_/Y _13693_/X VGND VGND VPWR VPWR _13732_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__25475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_40_0_HCLK clkbuf_5_20_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16451_ _19091_/A VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__buf_2
XFILLER_232_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13663_ _13662_/X VGND VGND VPWR VPWR _13664_/B sky130_fd_sc_hd__inv_2
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15402_ _15411_/A _15401_/X VGND VGND VPWR VPWR _15409_/B sky130_fd_sc_hd__or2_4
X_12614_ _12710_/B VGND VGND VPWR VPWR _12702_/A sky130_fd_sc_hd__buf_2
X_19170_ _19165_/Y _19168_/X _19169_/X _19168_/X VGND VGND VPWR VPWR _19170_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16382_ _16382_/A _16382_/B VGND VGND VPWR VPWR _16390_/A sky130_fd_sc_hd__nor2_4
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22666__A1 _15718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13594_ _25261_/Q _13561_/Y _13857_/A _14569_/B VGND VGND VPWR VPWR _13594_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22666__B2 _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18121_ _18084_/X _23904_/Q VGND VGND VPWR VPWR _18122_/C sky130_fd_sc_hd__or2_4
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15333_ _15355_/A _15331_/X _15332_/X VGND VGND VPWR VPWR _25010_/D sky130_fd_sc_hd__and3_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12545_ _12545_/A VGND VGND VPWR VPWR _12545_/Y sky130_fd_sc_hd__inv_2
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18052_ _18090_/A _23890_/Q VGND VGND VPWR VPWR _18052_/X sky130_fd_sc_hd__or2_4
XFILLER_200_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15264_ _15255_/X _15262_/X _15264_/C VGND VGND VPWR VPWR _15264_/X sky130_fd_sc_hd__and3_4
XFILLER_185_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12476_ _12514_/A VGND VGND VPWR VPWR _12501_/A sky130_fd_sc_hd__buf_2
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17003_ _17159_/A VGND VGND VPWR VPWR _17139_/A sky130_fd_sc_hd__inv_2
X_14215_ _20525_/A _14208_/X _13849_/X _14210_/X VGND VGND VPWR VPWR _14215_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22969__A2 _22851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ _15195_/A _15195_/B VGND VGND VPWR VPWR _15197_/B sky130_fd_sc_hd__or2_4
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14146_ _14119_/X _14144_/X _14430_/A _14145_/X VGND VGND VPWR VPWR _14146_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__17845__A1 _17766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14077_ _14021_/B _14074_/X _14066_/X _14058_/C _14075_/X VGND VGND VPWR VPWR _14077_/X
+ sky130_fd_sc_hd__a32o_4
X_18954_ _23918_/Q VGND VGND VPWR VPWR _18954_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21929__B1 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13028_ _13027_/X VGND VGND VPWR VPWR _13028_/Y sky130_fd_sc_hd__inv_2
X_17905_ _22005_/A _17904_/X VGND VGND VPWR VPWR _17905_/Y sky130_fd_sc_hd__nand2_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18885_ _23958_/Q _18885_/B VGND VGND VPWR VPWR _18886_/B sky130_fd_sc_hd__or2_4
XFILLER_239_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17836_ _16933_/A _17836_/B VGND VGND VPWR VPWR _17836_/X sky130_fd_sc_hd__or2_4
XFILLER_239_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_245_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17767_ _17767_/A VGND VGND VPWR VPWR _17768_/D sky130_fd_sc_hd__inv_2
X_14979_ _14910_/Y _24445_/Q _25033_/Q _14978_/Y VGND VGND VPWR VPWR _14983_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19506_ _19965_/A _18285_/D _19505_/X VGND VGND VPWR VPWR _19507_/A sky130_fd_sc_hd__or3_4
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16718_ _24488_/Q VGND VGND VPWR VPWR _16718_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17698_ _17537_/Y _17671_/X VGND VGND VPWR VPWR _17703_/B sky130_fd_sc_hd__or2_4
XFILLER_222_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19437_ _19436_/X VGND VGND VPWR VPWR _19438_/A sky130_fd_sc_hd__inv_2
X_16649_ _15565_/X _15651_/X VGND VGND VPWR VPWR _16652_/A sky130_fd_sc_hd__or2_4
XFILLER_211_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19368_ _19368_/A VGND VGND VPWR VPWR _19368_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18319_ _18319_/A VGND VGND VPWR VPWR _21463_/A sky130_fd_sc_hd__inv_2
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19299_ _23796_/Q VGND VGND VPWR VPWR _19299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12517__A _21083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21330_ _21330_/A VGND VGND VPWR VPWR _21330_/X sky130_fd_sc_hd__buf_2
XFILLER_163_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_60_0_HCLK clkbuf_8_61_0_HCLK/A VGND VGND VPWR VPWR _24952_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_190_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21261_ _21255_/X _21260_/X _14692_/A VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__o21a_4
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24780__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21549__B _21719_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23000_ _17322_/A _22926_/X _12857_/A _22927_/X VGND VGND VPWR VPWR _23000_/X sky130_fd_sc_hd__a2bb2o_4
X_20212_ _13757_/C _13761_/X _13744_/X _13770_/X VGND VGND VPWR VPWR _20213_/A sky130_fd_sc_hd__or4_4
X_21192_ _21211_/A _21192_/B VGND VGND VPWR VPWR _21193_/C sky130_fd_sc_hd__or2_4
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24960__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15847__B1 _15486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20143_ _23502_/Q VGND VGND VPWR VPWR _21403_/B sky130_fd_sc_hd__inv_2
XANTENNA__20840__B1 _20836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19038__B1 _19012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20074_ _23526_/Q VGND VGND VPWR VPWR _20074_/Y sky130_fd_sc_hd__inv_2
X_24951_ _25103_/CLK _15505_/X HRESETn VGND VGND VPWR VPWR _17456_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21565__A _21565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23902_ _25082_/CLK _23902_/D VGND VGND VPWR VPWR _18996_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_246_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24882_ _24889_/CLK _15740_/X HRESETn VGND VGND VPWR VPWR _12595_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16272__B1 _15483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23833_ _24100_/CLK _23833_/D VGND VGND VPWR VPWR _23833_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23764_ _25077_/CLK _19393_/X VGND VGND VPWR VPWR _17956_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _20976_/A _13529_/A VGND VGND VPWR VPWR _24108_/D sky130_fd_sc_hd__and2_4
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25503_ _25177_/CLK _11991_/X HRESETn VGND VGND VPWR VPWR _11663_/C sky130_fd_sc_hd__dfrtp_4
Xclkbuf_5_27_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22715_ _21879_/A _22715_/B _22714_/X VGND VGND VPWR VPWR _22715_/X sky130_fd_sc_hd__and3_4
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23695_ _23717_/CLK _19588_/X VGND VGND VPWR VPWR _19586_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25434_ _25419_/CLK _12650_/Y HRESETn VGND VGND VPWR VPWR _25434_/Q sky130_fd_sc_hd__dfrtp_4
X_22646_ _24629_/Q _22610_/B VGND VGND VPWR VPWR _22646_/X sky130_fd_sc_hd__or2_4
XFILLER_186_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25365_ _25365_/CLK _13042_/X HRESETn VGND VGND VPWR VPWR _25365_/Q sky130_fd_sc_hd__dfrtp_4
X_22577_ _22577_/A _22577_/B VGND VGND VPWR VPWR _22577_/X sky130_fd_sc_hd__and2_4
XANTENNA__24868__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12330_ _24849_/Q VGND VGND VPWR VPWR _12330_/Y sky130_fd_sc_hd__inv_2
X_24316_ _25543_/CLK _24316_/D HRESETn VGND VGND VPWR VPWR _24316_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21528_ _21326_/X _21425_/X _21528_/C _21527_/X VGND VGND VPWR VPWR HRDATA[1] sky130_fd_sc_hd__or4_4
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25296_ _24378_/CLK _25296_/D HRESETn VGND VGND VPWR VPWR _11688_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21871__A2 _22424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ _25460_/Q VGND VGND VPWR VPWR _12261_/Y sky130_fd_sc_hd__inv_2
X_24247_ _23754_/CLK _24247_/D HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15738__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21459_ _16936_/X _21457_/X _12513_/A _22447_/A VGND VGND VPWR VPWR _21459_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23073__B2 _21229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14000_ _25246_/Q _25245_/Q _14000_/C VGND VGND VPWR VPWR _14021_/D sky130_fd_sc_hd__or3_4
XFILLER_135_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _25444_/Q _12190_/Y _12191_/Y _23196_/A VGND VGND VPWR VPWR _12192_/X sky130_fd_sc_hd__a2bb2o_4
X_24178_ _23973_/CLK _18553_/X HRESETn VGND VGND VPWR VPWR _24178_/Q sky130_fd_sc_hd__dfrtp_4
X_23129_ _15553_/X VGND VGND VPWR VPWR _23129_/X sky130_fd_sc_hd__buf_2
XFILLER_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15951_ _12264_/Y _15947_/X _15950_/X _15947_/X VGND VGND VPWR VPWR _15951_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15853__A3 _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14902_ _14902_/A VGND VGND VPWR VPWR _14902_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15882_ _15858_/X _15865_/X _15732_/X _23162_/A _15872_/X VGND VGND VPWR VPWR _24816_/D
+ sky130_fd_sc_hd__a32o_4
X_18670_ _18670_/A VGND VGND VPWR VPWR _18717_/A sky130_fd_sc_hd__buf_2
XFILLER_237_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17621_ _17663_/A _17590_/X _17553_/Y _17621_/D VGND VGND VPWR VPWR _17621_/X sky130_fd_sc_hd__or4_4
X_14833_ _14832_/X VGND VGND VPWR VPWR _14852_/A sky130_fd_sc_hd__buf_2
XANTENNA__24001__D scl_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ _21240_/A VGND VGND VPWR VPWR _21248_/A sky130_fd_sc_hd__inv_2
X_17552_ _11768_/Y _24322_/Q _25545_/Q _17579_/B VGND VGND VPWR VPWR _17552_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19201__B1 _19131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17510__A1_N _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11976_ _11970_/C _11970_/D _11713_/Y _25505_/Q VGND VGND VPWR VPWR _11976_/X sky130_fd_sc_hd__and4_4
XFILLER_245_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22887__B2 _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19599__B _13782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16015__B1 _15950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13715_ _13711_/B _13689_/X _13714_/X _13712_/X _13702_/A VGND VGND VPWR VPWR _25298_/D
+ sky130_fd_sc_hd__a32o_4
X_16503_ _16502_/Y _16500_/X _16417_/X _16500_/X VGND VGND VPWR VPWR _24570_/D sky130_fd_sc_hd__a2bb2o_4
X_17483_ _18938_/B _17474_/X _17481_/Y _17482_/Y VGND VGND VPWR VPWR _17484_/D sky130_fd_sc_hd__a211o_4
X_14695_ _14706_/A _14695_/B VGND VGND VPWR VPWR _14695_/Y sky130_fd_sc_hd__nor2_4
XFILLER_189_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19222_ _18136_/B VGND VGND VPWR VPWR _19222_/Y sky130_fd_sc_hd__inv_2
X_13646_ _13645_/X VGND VGND VPWR VPWR _13647_/A sky130_fd_sc_hd__inv_2
X_16434_ _16434_/A VGND VGND VPWR VPWR _16434_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _16290_/A VGND VGND VPWR VPWR _16365_/X sky130_fd_sc_hd__buf_2
X_19153_ _19150_/Y _19145_/X _19151_/X _19152_/X VGND VGND VPWR VPWR _19153_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A VGND VGND VPWR VPWR _14586_/C sky130_fd_sc_hd__buf_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15316_ _15346_/A _15345_/C _15303_/X _15315_/X VGND VGND VPWR VPWR _15316_/X sky130_fd_sc_hd__or4_4
X_18104_ _18168_/A _18104_/B VGND VGND VPWR VPWR _18104_/X sky130_fd_sc_hd__or2_4
XFILLER_185_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12528_ _12520_/X _12522_/X _12525_/X _12527_/X VGND VGND VPWR VPWR _12567_/A sky130_fd_sc_hd__or4_4
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16296_ _16296_/A VGND VGND VPWR VPWR _16296_/Y sky130_fd_sc_hd__inv_2
X_19084_ _13307_/B VGND VGND VPWR VPWR _19084_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21862__A2 _22176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_47_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15247_ _15073_/X _15294_/A VGND VGND VPWR VPWR _15247_/X sky130_fd_sc_hd__or2_4
X_18035_ _17985_/A VGND VGND VPWR VPWR _18036_/A sky130_fd_sc_hd__buf_2
XFILLER_172_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12459_ _12197_/X _12449_/D _12411_/X _12457_/B VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18024__A _18013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15178_ _15178_/A _15176_/A VGND VGND VPWR VPWR _15178_/X sky130_fd_sc_hd__or2_4
XANTENNA__20417__A3 _14248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23947__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15829__B1 _24840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14129_ _14114_/Y _14128_/X VGND VGND VPWR VPWR _14129_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19986_ _17733_/A VGND VGND VPWR VPWR _19986_/X sky130_fd_sc_hd__buf_2
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _17477_/A _18937_/B _18333_/C VGND VGND VPWR VPWR _18938_/C sky130_fd_sc_hd__or3_4
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19440__B1 _19439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ _16466_/Y _18606_/X _16466_/Y _18606_/X VGND VGND VPWR VPWR _18868_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17819_ _17766_/A _17766_/B _17818_/X VGND VGND VPWR VPWR _17820_/B sky130_fd_sc_hd__or3_4
XFILLER_243_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18799_ _18805_/A _18799_/B _18799_/C VGND VGND VPWR VPWR _18799_/X sky130_fd_sc_hd__or3_4
X_20830_ _20830_/A VGND VGND VPWR VPWR _20831_/A sky130_fd_sc_hd__inv_2
XFILLER_70_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20761_ _20788_/A VGND VGND VPWR VPWR _20761_/X sky130_fd_sc_hd__buf_2
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22500_ _22500_/A VGND VGND VPWR VPWR _22500_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23480_ _23488_/CLK _23480_/D VGND VGND VPWR VPWR _23480_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692_ _23386_/D VGND VGND VPWR VPWR _20693_/A sky130_fd_sc_hd__inv_2
XFILLER_195_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22944__A _22944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22431_ _21034_/X VGND VGND VPWR VPWR _22431_/X sky130_fd_sc_hd__buf_2
XFILLER_176_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25150_ _25223_/CLK _14421_/X HRESETn VGND VGND VPWR VPWR _14414_/A sky130_fd_sc_hd__dfstp_4
X_22362_ _22036_/A _22362_/B _22362_/C VGND VGND VPWR VPWR _22362_/X sky130_fd_sc_hd__and3_4
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24101_ _24101_/CLK _20969_/X HRESETn VGND VGND VPWR VPWR RsTx_S1 sky130_fd_sc_hd__dfstp_4
XFILLER_163_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21313_ _21300_/Y VGND VGND VPWR VPWR _21314_/A sky130_fd_sc_hd__buf_2
XFILLER_136_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25081_ _25082_/CLK _25081_/D HRESETn VGND VGND VPWR VPWR _13613_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22293_ _21082_/X _22287_/X _22836_/A _22292_/X VGND VGND VPWR VPWR _22294_/B sky130_fd_sc_hd__a22oi_4
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24032_ _24495_/CLK _24032_/D HRESETn VGND VGND VPWR VPWR _20776_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17809__A1 _17753_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21244_ _21275_/A _21244_/B _21243_/X VGND VGND VPWR VPWR _21244_/X sky130_fd_sc_hd__and3_4
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_4_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21175_ _21874_/A _21175_/B _21174_/X VGND VGND VPWR VPWR _21175_/X sky130_fd_sc_hd__and3_4
XANTENNA__16493__B1 _16407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20126_ _20126_/A VGND VGND VPWR VPWR _22382_/B sky130_fd_sc_hd__inv_2
XFILLER_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16389__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15293__A _15293_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _23532_/Q VGND VGND VPWR VPWR _20057_/Y sky130_fd_sc_hd__inv_2
X_24934_ _25093_/CLK _15545_/X HRESETn VGND VGND VPWR VPWR _11731_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_245_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20289__A2_N _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24865_ _24476_/CLK _15773_/X HRESETn VGND VGND VPWR VPWR _12572_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22318__B1 _15676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ HWDATA[10] VGND VGND VPWR VPWR _11830_/X sky130_fd_sc_hd__buf_2
X_23816_ _23454_/CLK _19247_/X VGND VGND VPWR VPWR _13349_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24796_ _24799_/CLK _15911_/X HRESETn VGND VGND VPWR VPWR _22302_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23015__A _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11757_/Y _11751_/X _11758_/X _11760_/X VGND VGND VPWR VPWR _25554_/D sky130_fd_sc_hd__a2bb2o_4
X_23747_ _23669_/CLK _23747_/D VGND VGND VPWR VPWR _17995_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20836_/X _20958_/Y _16659_/A _20883_/A VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18870__A1_N _16482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _25323_/Q VGND VGND VPWR VPWR _13500_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14477_/Y _14475_/X _14479_/X _14475_/X VGND VGND VPWR VPWR _25128_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _24232_/Q VGND VGND VPWR VPWR _11692_/Y sky130_fd_sc_hd__inv_2
X_23678_ _23678_/CLK _19647_/X VGND VGND VPWR VPWR _19645_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13315_/A _13427_/X _13430_/X VGND VGND VPWR VPWR _13431_/X sky130_fd_sc_hd__or3_4
X_25417_ _25419_/CLK _12720_/X HRESETn VGND VGND VPWR VPWR _12519_/A sky130_fd_sc_hd__dfrtp_4
X_22629_ _22592_/A _22629_/B _22628_/X VGND VGND VPWR VPWR _22629_/X sky130_fd_sc_hd__and3_4
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20227__A2_N _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16150_ _22574_/A VGND VGND VPWR VPWR _16150_/Y sky130_fd_sc_hd__inv_2
X_13362_ _13245_/X _13362_/B VGND VGND VPWR VPWR _13363_/C sky130_fd_sc_hd__or2_4
X_25348_ _25358_/CLK _25348_/D HRESETn VGND VGND VPWR VPWR _25348_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24631__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15101_ _15101_/A VGND VGND VPWR VPWR _15396_/A sky130_fd_sc_hd__inv_2
X_12313_ _12312_/X _24841_/Q _12311_/Y _24841_/Q VGND VGND VPWR VPWR _12322_/A sky130_fd_sc_hd__a2bb2o_4
X_16081_ _16080_/Y _16076_/X _15995_/X _16076_/X VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__a2bb2o_4
X_13293_ _13290_/X _13293_/B _13292_/X VGND VGND VPWR VPWR _13293_/X sky130_fd_sc_hd__and3_4
X_25279_ _23647_/CLK _13810_/X HRESETn VGND VGND VPWR VPWR _25279_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15032_ _15032_/A VGND VGND VPWR VPWR _15032_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21057__B1 _21882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12244_ _12296_/B VGND VGND VPWR VPWR _12439_/B sky130_fd_sc_hd__buf_2
XFILLER_6_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18779__A _18710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19840_ _22371_/B _19839_/X _19790_/X _19839_/X VGND VGND VPWR VPWR _23612_/D sky130_fd_sc_hd__a2bb2o_4
X_12175_ _12175_/A _25172_/Q VGND VGND VPWR VPWR _12175_/X sky130_fd_sc_hd__and2_4
XANTENNA__19670__B1 _19454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16484__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19771_ _13299_/B VGND VGND VPWR VPWR _19771_/Y sky130_fd_sc_hd__inv_2
X_16983_ _24386_/Q VGND VGND VPWR VPWR _17142_/A sky130_fd_sc_hd__inv_2
XFILLER_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18722_ _18717_/A _18711_/X _18714_/X _18719_/B VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__a211o_4
XFILLER_209_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15934_ _15668_/B _15934_/B VGND VGND VPWR VPWR _15934_/X sky130_fd_sc_hd__or2_4
XFILLER_237_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16236__B1 _11805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18653_ _16599_/Y _18782_/A _16599_/Y _18782_/A VGND VGND VPWR VPWR _18659_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22572__A3 _21550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15865_ _15895_/A VGND VGND VPWR VPWR _15865_/X sky130_fd_sc_hd__buf_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22309__B1 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17604_ _17569_/X _17616_/B VGND VGND VPWR VPWR _17604_/X sky130_fd_sc_hd__or2_4
X_14816_ _14816_/A _14816_/B _14816_/C VGND VGND VPWR VPWR _14817_/A sky130_fd_sc_hd__or3_4
X_18584_ _18400_/Y _18568_/X VGND VGND VPWR VPWR _18586_/B sky130_fd_sc_hd__nand2_4
X_15796_ _15844_/A VGND VGND VPWR VPWR _15796_/X sky130_fd_sc_hd__buf_2
XFILLER_240_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17535_ _17535_/A VGND VGND VPWR VPWR _17578_/B sky130_fd_sc_hd__inv_2
X_11959_ _20010_/A VGND VGND VPWR VPWR _19646_/A sky130_fd_sc_hd__buf_2
X_14747_ _14735_/X _14739_/Y VGND VGND VPWR VPWR _14747_/Y sky130_fd_sc_hd__nor2_4
XFILLER_199_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13451__A _13451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14678_ _13626_/A VGND VGND VPWR VPWR _19166_/A sky130_fd_sc_hd__buf_2
X_17466_ _17466_/A VGND VGND VPWR VPWR _18347_/A sky130_fd_sc_hd__inv_2
XANTENNA__24719__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19205_ _19205_/A VGND VGND VPWR VPWR _19205_/Y sky130_fd_sc_hd__inv_2
X_13629_ _13628_/X VGND VGND VPWR VPWR _14670_/A sky130_fd_sc_hd__inv_2
X_16417_ HWDATA[18] VGND VGND VPWR VPWR _16417_/X sky130_fd_sc_hd__buf_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17397_ _20627_/A _20624_/A VGND VGND VPWR VPWR _17398_/B sky130_fd_sc_hd__or2_4
XANTENNA__16762__A _16762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19136_ _13411_/B VGND VGND VPWR VPWR _19136_/Y sky130_fd_sc_hd__inv_2
X_16348_ _16348_/A VGND VGND VPWR VPWR _16348_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11784__B1 _11783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16279_ _16278_/Y _16196_/X _15489_/X _16196_/X VGND VGND VPWR VPWR _24652_/D sky130_fd_sc_hd__a2bb2o_4
X_19067_ _19067_/A VGND VGND VPWR VPWR _19067_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18018_ _18098_/A VGND VGND VPWR VPWR _18060_/A sky130_fd_sc_hd__buf_2
XFILLER_172_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14722__B1 _14721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_134_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23669_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_197_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24493_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19969_ _23563_/Q VGND VGND VPWR VPWR _19969_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22004__A _22003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22980_ _21101_/X VGND VGND VPWR VPWR _23208_/A sky130_fd_sc_hd__buf_2
XFILLER_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21931_ _17727_/A _21931_/B VGND VGND VPWR VPWR _21931_/X sky130_fd_sc_hd__or2_4
X_24650_ _24651_/CLK _24650_/D HRESETn VGND VGND VPWR VPWR _24650_/Q sky130_fd_sc_hd__dfrtp_4
X_21862_ _20514_/D _22176_/B _14470_/Y _17424_/X VGND VGND VPWR VPWR _21863_/D sky130_fd_sc_hd__o22a_4
XFILLER_36_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23601_ _23488_/CLK _23601_/D VGND VGND VPWR VPWR _23601_/Q sky130_fd_sc_hd__dfxtp_4
X_20813_ _13145_/X VGND VGND VPWR VPWR _20818_/B sky130_fd_sc_hd__inv_2
XANTENNA__15560__B _21122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19716__B2 _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24581_ _24562_/CLK _16477_/X HRESETn VGND VGND VPWR VPWR _16474_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21793_ _21789_/X _21792_/X _14758_/X VGND VGND VPWR VPWR _21793_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21523__A1 _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23514_/CLK _23532_/D VGND VGND VPWR VPWR _23532_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20744_ _20744_/A VGND VGND VPWR VPWR _20744_/X sky130_fd_sc_hd__buf_2
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ _23466_/CLK _20250_/X VGND VGND VPWR VPWR _20247_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20675_ _20675_/A _20675_/B _20675_/C VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__and3_4
XFILLER_149_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16688__A1_N _16687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16672__A _16653_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25202_ _25204_/CLK _14243_/X HRESETn VGND VGND VPWR VPWR _25202_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ _23027_/B _22413_/X _22303_/X VGND VGND VPWR VPWR _22414_/X sky130_fd_sc_hd__and3_4
X_23394_ _23522_/CLK _23394_/D VGND VGND VPWR VPWR _20422_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_195_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25133_ _25137_/CLK _25133_/D HRESETn VGND VGND VPWR VPWR _14465_/A sky130_fd_sc_hd__dfrtp_4
X_22345_ _21949_/A _22343_/X _22344_/X VGND VGND VPWR VPWR _22345_/X sky130_fd_sc_hd__and3_4
XANTENNA__24042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16611__A1_N _16608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_30_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_25064_ _24258_/CLK _25064_/D HRESETn VGND VGND VPWR VPWR _14783_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22276_ _23402_/Q _22013_/Y _22524_/B _22275_/X VGND VGND VPWR VPWR _22277_/A sky130_fd_sc_hd__a211o_4
XFILLER_191_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_93_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24015_ _24015_/CLK _20700_/Y HRESETn VGND VGND VPWR VPWR _13131_/B sky130_fd_sc_hd__dfrtp_4
X_21227_ _24047_/Q VGND VGND VPWR VPWR _21227_/Y sky130_fd_sc_hd__inv_2
X_21158_ _20548_/B VGND VGND VPWR VPWR _21158_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16626__A1_N _16625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20109_ _20100_/Y VGND VGND VPWR VPWR _20109_/X sky130_fd_sc_hd__buf_2
XFILLER_219_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13980_ _13980_/A VGND VGND VPWR VPWR _13980_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21089_ _15866_/X VGND VGND VPWR VPWR _21090_/A sky130_fd_sc_hd__buf_2
XANTENNA__16218__B1 _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12931_ _12921_/C _12921_/D _12883_/X _12929_/B VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__a211o_4
XFILLER_207_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24917_ _24825_/CLK _15600_/X HRESETn VGND VGND VPWR VPWR _15599_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22568__B _21450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12862_ _12817_/Y _12825_/Y _12862_/C _12895_/B VGND VGND VPWR VPWR _12862_/X sky130_fd_sc_hd__or4_4
X_15650_ _22121_/A VGND VGND VPWR VPWR _15650_/X sky130_fd_sc_hd__buf_2
X_24848_ _24878_/CLK _15816_/X HRESETn VGND VGND VPWR VPWR _24848_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _16241_/A VGND VGND VPWR VPWR _11813_/X sky130_fd_sc_hd__buf_2
X_14601_ _14601_/A _14577_/B VGND VGND VPWR VPWR _14601_/Y sky130_fd_sc_hd__nand2_4
XFILLER_215_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15581_/A VGND VGND VPWR VPWR _15581_/Y sky130_fd_sc_hd__inv_2
X_12793_ _12793_/A VGND VGND VPWR VPWR _12855_/A sky130_fd_sc_hd__inv_2
X_24779_ _24803_/CLK _15955_/X HRESETn VGND VGND VPWR VPWR _24779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24883__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15992__A2 _15895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14530_/X _14531_/X _25124_/Q _14526_/X VGND VGND VPWR VPWR _25112_/D sky130_fd_sc_hd__o22a_4
X_17320_ _17322_/B VGND VGND VPWR VPWR _17321_/B sky130_fd_sc_hd__inv_2
XANTENNA__22456__A1_N _17364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _21332_/A VGND VGND VPWR VPWR _11744_/X sky130_fd_sc_hd__buf_2
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24812__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20166__A2_N _20163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14468_/A VGND VGND VPWR VPWR _14463_/X sky130_fd_sc_hd__buf_2
X_17251_ _17251_/A VGND VGND VPWR VPWR _17252_/D sky130_fd_sc_hd__inv_2
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11675_/A _11675_/B _11675_/C _11674_/X VGND VGND VPWR VPWR _11709_/A sky130_fd_sc_hd__or4_4
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13317_/A _13414_/B VGND VGND VPWR VPWR _13415_/C sky130_fd_sc_hd__or2_4
X_16202_ _16202_/A VGND VGND VPWR VPWR _16227_/A sky130_fd_sc_hd__buf_2
XFILLER_169_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _16331_/Y _17262_/A _16331_/Y _17262_/A VGND VGND VPWR VPWR _17190_/A sky130_fd_sc_hd__a2bb2o_4
X_14394_ _20463_/A _14391_/X _13844_/X _14393_/X VGND VGND VPWR VPWR _25158_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15820__A1_N _12375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16133_ _16132_/Y _16128_/X _15972_/X _16128_/X VGND VGND VPWR VPWR _16133_/X sky130_fd_sc_hd__a2bb2o_4
X_13345_ _13212_/A VGND VGND VPWR VPWR _13410_/A sky130_fd_sc_hd__buf_2
XFILLER_127_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16064_ _16063_/Y _16061_/X _15767_/X _16061_/X VGND VGND VPWR VPWR _24729_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14704__B1 _21630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13276_ _13217_/X _13274_/X _13275_/X VGND VGND VPWR VPWR _13276_/X sky130_fd_sc_hd__and3_4
XFILLER_170_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15015_ _15188_/A _24480_/Q _15182_/A _15014_/Y VGND VGND VPWR VPWR _15021_/B sky130_fd_sc_hd__o22a_4
X_12227_ _25467_/Q _24782_/Q _12225_/Y _12226_/Y VGND VGND VPWR VPWR _12235_/B sky130_fd_sc_hd__o22a_4
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_207_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _24528_/CLK sky130_fd_sc_hd__clkbuf_1
X_19823_ _19821_/Y _19816_/X _19772_/X _19822_/X VGND VGND VPWR VPWR _23618_/D sky130_fd_sc_hd__a2bb2o_4
X_12158_ _24118_/Q _12138_/A _12157_/Y VGND VGND VPWR VPWR _12158_/X sky130_fd_sc_hd__o21a_4
XFILLER_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ _19752_/Y _19748_/X _19753_/X _19748_/X VGND VGND VPWR VPWR _23640_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12089_ _12087_/Y _12083_/X _11851_/X _12088_/X VGND VGND VPWR VPWR _12089_/X sky130_fd_sc_hd__a2bb2o_4
X_16966_ _21022_/B _16964_/X _16965_/Y VGND VGND VPWR VPWR _24410_/D sky130_fd_sc_hd__o21a_4
XFILLER_238_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18705_ _18720_/A _18717_/A _18678_/Y _18717_/B VGND VGND VPWR VPWR _18705_/X sky130_fd_sc_hd__or4_4
XANTENNA__21663__A _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15917_ _12804_/Y _15912_/X _15848_/X _15880_/A VGND VGND VPWR VPWR _15917_/X sky130_fd_sc_hd__a2bb2o_4
X_19685_ _19684_/Y _19682_/X _19560_/X _19682_/X VGND VGND VPWR VPWR _19685_/X sky130_fd_sc_hd__a2bb2o_4
X_16897_ _19810_/A VGND VGND VPWR VPWR _16897_/X sky130_fd_sc_hd__buf_2
XFILLER_209_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21753__A1 _16625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18636_ _16558_/A _24160_/Q _16558_/Y _18720_/A VGND VGND VPWR VPWR _18636_/X sky130_fd_sc_hd__o22a_4
X_15848_ _14479_/A VGND VGND VPWR VPWR _15848_/X sky130_fd_sc_hd__buf_2
XFILLER_224_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18567_ _18480_/Y _18566_/X VGND VGND VPWR VPWR _18567_/X sky130_fd_sc_hd__or2_4
XFILLER_224_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15779_ _12561_/Y _15772_/X _15486_/X _15772_/X VGND VGND VPWR VPWR _24862_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17518_ _24304_/Q VGND VGND VPWR VPWR _17518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24553__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18498_ _18488_/C _18510_/B VGND VGND VPWR VPWR _18499_/A sky130_fd_sc_hd__or2_4
XFILLER_21_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22494__A _22721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17449_ _17448_/X VGND VGND VPWR VPWR _17450_/B sky130_fd_sc_hd__buf_2
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20460_ _20460_/A VGND VGND VPWR VPWR _20461_/D sky130_fd_sc_hd__inv_2
XFILLER_220_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ _18938_/A _19075_/B _19119_/C VGND VGND VPWR VPWR _19119_/X sky130_fd_sc_hd__or3_4
X_20391_ _20385_/Y VGND VGND VPWR VPWR _20391_/X sky130_fd_sc_hd__buf_2
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22130_ _15476_/Y _21370_/X _14237_/Y _14230_/A VGND VGND VPWR VPWR _22131_/A sky130_fd_sc_hd__o22a_4
XFILLER_133_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_133_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21838__A _13793_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22769__B1 _21844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22061_ _22058_/Y _22059_/X _21981_/X _22060_/X VGND VGND VPWR VPWR _23354_/B sky130_fd_sc_hd__a211o_4
XANTENNA__19308__A _19151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18212__A _18051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21012_ _23984_/Q VGND VGND VPWR VPWR _21012_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13356__A _13356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21992__B2 _20356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22963_ _20923_/Y _22842_/X _20785_/A _22298_/A VGND VGND VPWR VPWR _22963_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16667__A _16654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21914_ _21914_/A _20179_/Y VGND VGND VPWR VPWR _21916_/B sky130_fd_sc_hd__or2_4
X_24702_ _24756_/CLK _24702_/D HRESETn VGND VGND VPWR VPWR _22792_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15571__A _15626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22894_ _20775_/Y _21124_/X _20914_/Y _21229_/X VGND VGND VPWR VPWR _22894_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24633_ _24629_/CLK _24633_/D HRESETn VGND VGND VPWR VPWR _24633_/Q sky130_fd_sc_hd__dfrtp_4
X_21845_ _22947_/A VGND VGND VPWR VPWR _22695_/B sky130_fd_sc_hd__buf_2
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24564_ _24566_/CLK _24564_/D HRESETn VGND VGND VPWR VPWR _16517_/A sky130_fd_sc_hd__dfrtp_4
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ _21772_/X _21775_/X _14758_/X VGND VGND VPWR VPWR _21776_/X sky130_fd_sc_hd__o21a_4
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23516_/CLK _20106_/X VGND VGND VPWR VPWR _23515_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20727_ _20725_/A _20725_/B _20731_/B VGND VGND VPWR VPWR _20727_/Y sky130_fd_sc_hd__a21oi_4
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24495_ _24495_/CLK _24495_/D HRESETn VGND VGND VPWR VPWR _16701_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _23926_/CLK _23446_/D VGND VGND VPWR VPWR _23446_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20658_ _14247_/Y _20646_/X _20637_/X _20657_/X VGND VGND VPWR VPWR _20659_/A sky130_fd_sc_hd__a211o_4
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23377_ _21020_/X VGND VGND VPWR VPWR IRQ[21] sky130_fd_sc_hd__buf_2
X_20589_ _18885_/B _20588_/Y _20597_/C VGND VGND VPWR VPWR _20589_/X sky130_fd_sc_hd__and3_4
XFILLER_180_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13130_ _24017_/Q VGND VGND VPWR VPWR _13130_/Y sky130_fd_sc_hd__inv_2
X_25116_ _24095_/CLK _14518_/X HRESETn VGND VGND VPWR VPWR _25116_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18140__A3 _18139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22328_ _17198_/X _21321_/A _12218_/A _21081_/A VGND VGND VPWR VPWR _22328_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13061_ _12997_/D _13061_/B VGND VGND VPWR VPWR _13074_/A sky130_fd_sc_hd__or2_4
X_25047_ _25212_/CLK _14888_/Y HRESETn VGND VGND VPWR VPWR _14873_/B sky130_fd_sc_hd__dfrtp_4
X_22259_ _21679_/A _22251_/X _22258_/X VGND VGND VPWR VPWR _22259_/X sky130_fd_sc_hd__and3_4
XFILLER_140_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23385__D scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ _25315_/Q _20971_/A _25315_/Q _20971_/A VGND VGND VPWR VPWR _12012_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16439__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25082__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21983__A1 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16820_ _16810_/X VGND VGND VPWR VPWR _16820_/X sky130_fd_sc_hd__buf_2
XANTENNA__25011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_180_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _23954_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_37_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _23494_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21483__A _21675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16751_ _16750_/Y _16748_/X _15734_/X _16748_/X VGND VGND VPWR VPWR _16751_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13963_ _13963_/A _13963_/B _13955_/A _13913_/Y VGND VGND VPWR VPWR _13963_/X sky130_fd_sc_hd__or4_4
X_15702_ _18029_/A VGND VGND VPWR VPWR _15703_/A sky130_fd_sc_hd__inv_2
XFILLER_206_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12914_ _12834_/Y _12913_/X VGND VGND VPWR VPWR _12917_/B sky130_fd_sc_hd__or2_4
X_19470_ _19470_/A VGND VGND VPWR VPWR _19470_/Y sky130_fd_sc_hd__inv_2
X_13894_ _13893_/X VGND VGND VPWR VPWR _13982_/A sky130_fd_sc_hd__buf_2
X_16682_ _16682_/A VGND VGND VPWR VPWR _16682_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18421_ _24192_/Q VGND VGND VPWR VPWR _18488_/B sky130_fd_sc_hd__inv_2
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16611__B1 _16609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12845_ _12813_/X _12845_/B _12845_/C _12845_/D VGND VGND VPWR VPWR _12845_/X sky130_fd_sc_hd__or4_4
X_15633_ _15631_/Y _15626_/X _15632_/X _15626_/X VGND VGND VPWR VPWR _15633_/X sky130_fd_sc_hd__a2bb2o_4
X_18352_ _18352_/A VGND VGND VPWR VPWR _18352_/Y sky130_fd_sc_hd__inv_2
X_12776_ _25381_/Q VGND VGND VPWR VPWR _12777_/A sky130_fd_sc_hd__inv_2
X_15564_ _21172_/B VGND VGND VPWR VPWR _21855_/B sky130_fd_sc_hd__buf_2
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17305_/B VGND VGND VPWR VPWR _17303_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22160__B2 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A _12061_/B VGND VGND VPWR VPWR _15791_/D sky130_fd_sc_hd__or2_4
X_14515_ _23969_/Q VGND VGND VPWR VPWR _14515_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15493_/A _15493_/B _15494_/Y _14562_/Y VGND VGND VPWR VPWR _15495_/X sky130_fd_sc_hd__a211o_4
X_18283_ _17717_/X VGND VGND VPWR VPWR _18283_/X sky130_fd_sc_hd__buf_2
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _16367_/Y _17253_/A _24618_/Q _17391_/A VGND VGND VPWR VPWR _17238_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11658_/A VGND VGND VPWR VPWR _11661_/A sky130_fd_sc_hd__buf_2
X_14446_ _14446_/A VGND VGND VPWR VPWR _14446_/X sky130_fd_sc_hd__buf_2
XFILLER_174_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16518__A1_N _16517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _25161_/Q _14360_/A _25160_/Q _14354_/B VGND VGND VPWR VPWR _14377_/X sky130_fd_sc_hd__o22a_4
X_17165_ _17048_/Y _17166_/B VGND VGND VPWR VPWR _17165_/Y sky130_fd_sc_hd__nand2_4
XFILLER_128_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16462__D _15661_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22463__A2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16678__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ _13249_/A _23793_/Q VGND VGND VPWR VPWR _13330_/B sky130_fd_sc_hd__or2_4
X_16116_ _16103_/X VGND VGND VPWR VPWR _16116_/X sky130_fd_sc_hd__buf_2
XFILLER_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17096_ _17057_/D _17074_/X _17057_/B VGND VGND VPWR VPWR _17097_/C sky130_fd_sc_hd__o21a_4
XFILLER_115_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15656__A _13818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13259_ _13254_/X _13256_/X _13258_/X VGND VGND VPWR VPWR _13259_/X sky130_fd_sc_hd__and3_4
X_16047_ _16046_/Y _16044_/X _11809_/X _16044_/X VGND VGND VPWR VPWR _16047_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14560__A HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19806_ _19788_/Y VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__buf_2
X_17998_ _18006_/A VGND VGND VPWR VPWR _18189_/A sky130_fd_sc_hd__buf_2
XANTENNA__13607__C _25062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22489__A _23053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13113__C1 _13040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16850__B1 _16609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19737_ _19736_/Y _19733_/X _19692_/X _19733_/X VGND VGND VPWR VPWR _23646_/D sky130_fd_sc_hd__a2bb2o_4
X_16949_ _16166_/Y _24267_/Q _23237_/A _16957_/A VGND VGND VPWR VPWR _16954_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_244_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16487__A _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19668_ _19666_/Y _19667_/X _19566_/X _19667_/X VGND VGND VPWR VPWR _23671_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24734__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15405__A1 _15082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14208__A2 _14205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_8_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16602__B1 _16248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18619_ _24158_/Q VGND VGND VPWR VPWR _18703_/A sky130_fd_sc_hd__inv_2
XFILLER_92_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19599_ _13781_/A _13782_/A _19550_/C _19599_/D VGND VGND VPWR VPWR _19599_/X sky130_fd_sc_hd__and4_4
XANTENNA__22136__D1 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21630_ _21630_/A _21630_/B _21629_/X VGND VGND VPWR VPWR _21630_/X sky130_fd_sc_hd__and3_4
XFILLER_40_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23113__A _21126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21561_ _14434_/Y _14232_/A _14178_/Y _15471_/A VGND VGND VPWR VPWR _21563_/C sky130_fd_sc_hd__o22a_4
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18207__A _18013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16905__B2 _17767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23300_ _12275_/Y _21542_/X _24293_/Q _22501_/X VGND VGND VPWR VPWR _23302_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20512_ _20510_/X _20511_/X VGND VGND VPWR VPWR _20512_/X sky130_fd_sc_hd__or2_4
X_24280_ _24283_/CLK _17837_/X HRESETn VGND VGND VPWR VPWR _16933_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21492_ _21688_/A _21492_/B VGND VGND VPWR VPWR _21493_/C sky130_fd_sc_hd__or2_4
XFILLER_193_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23231_ _23231_/A _23119_/B VGND VGND VPWR VPWR _23231_/X sky130_fd_sc_hd__or2_4
X_20443_ _20445_/A _20443_/B VGND VGND VPWR VPWR _20443_/X sky130_fd_sc_hd__and2_4
XFILLER_193_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23162_ _23162_/A _23119_/B VGND VGND VPWR VPWR _23162_/X sky130_fd_sc_hd__or2_4
XFILLER_162_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20374_ _23415_/Q VGND VGND VPWR VPWR _20374_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22113_ _14450_/Y _14443_/A _14467_/Y _17424_/A VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19291__A2_N _19286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15566__A _15565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23093_ _23093_/A _23093_/B _23093_/C VGND VGND VPWR VPWR _23112_/B sky130_fd_sc_hd__and3_4
XANTENNA__19607__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25142__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22044_ _22040_/X _22043_/X _21697_/X VGND VGND VPWR VPWR _22044_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_253_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _24339_/CLK sky130_fd_sc_hd__clkbuf_1
X_23995_ _23998_/CLK _20663_/Y HRESETn VGND VGND VPWR VPWR _17404_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_216_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22946_ _24604_/Q _23189_/B VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__or2_4
XFILLER_56_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22877_ _23056_/A _22877_/B VGND VGND VPWR VPWR _22886_/C sky130_fd_sc_hd__and2_4
XANTENNA__18607__A1_N _16550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12630_ _12630_/A _12630_/B VGND VGND VPWR VPWR _12642_/D sky130_fd_sc_hd__or2_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ _21668_/A _21828_/B VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__or2_4
X_24616_ _25011_/CLK _24616_/D HRESETn VGND VGND VPWR VPWR _24616_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13562__A1_N _13560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12561_/A VGND VGND VPWR VPWR _12561_/Y sky130_fd_sc_hd__inv_2
X_24547_ _24542_/CLK _24547_/D HRESETn VGND VGND VPWR VPWR _16564_/A sky130_fd_sc_hd__dfrtp_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21759_ _21604_/A _21758_/X VGND VGND VPWR VPWR _21759_/Y sky130_fd_sc_hd__nor2_4
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14300_ _14300_/A _14305_/A _14303_/A _14303_/B VGND VGND VPWR VPWR _14300_/X sky130_fd_sc_hd__or4_4
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _15255_/X _15280_/B _15279_/Y VGND VGND VPWR VPWR _25019_/D sky130_fd_sc_hd__and3_4
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12229_/X _12489_/X VGND VGND VPWR VPWR _12493_/C sky130_fd_sc_hd__or2_4
X_24478_ _24473_/CLK _24478_/D HRESETn VGND VGND VPWR VPWR _24478_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _14204_/A VGND VGND VPWR VPWR _14232_/B sky130_fd_sc_hd__buf_2
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23429_ _23534_/CLK _23429_/D VGND VGND VPWR VPWR _20338_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15580__B1 _11766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22445__A2 _22444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24344__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14162_ _14124_/A _14124_/B _14124_/A _14124_/B VGND VGND VPWR VPWR _14162_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13113_ _13004_/B _13089_/X _13111_/B _13040_/X VGND VGND VPWR VPWR _13114_/A sky130_fd_sc_hd__a211o_4
X_14093_ _14068_/A VGND VGND VPWR VPWR _14093_/X sky130_fd_sc_hd__buf_2
X_18970_ _18968_/Y _18966_/X _18969_/X _18966_/X VGND VGND VPWR VPWR _23913_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_63_0_HCLK clkbuf_5_31_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _13044_/A _13044_/B _13043_/Y VGND VGND VPWR VPWR _13044_/X sky130_fd_sc_hd__and3_4
X_17921_ _24258_/Q VGND VGND VPWR VPWR _17921_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20208__B2 _20205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17691__A _17691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ _17852_/A _17850_/X _17851_/X VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__and3_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16803_ _16803_/A VGND VGND VPWR VPWR _16803_/Y sky130_fd_sc_hd__inv_2
X_17783_ _17775_/C _17782_/X _16964_/X _17776_/Y VGND VGND VPWR VPWR _17784_/A sky130_fd_sc_hd__a211o_4
X_14995_ _15067_/A VGND VGND VPWR VPWR _14996_/A sky130_fd_sc_hd__inv_2
XANTENNA__22102__A _15135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19522_ _19522_/A VGND VGND VPWR VPWR _21467_/B sky130_fd_sc_hd__inv_2
X_16734_ _16464_/A _16464_/B _22592_/A _21173_/C VGND VGND VPWR VPWR _16734_/X sky130_fd_sc_hd__and4_4
XFILLER_235_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13946_ _13964_/A VGND VGND VPWR VPWR _13958_/A sky130_fd_sc_hd__buf_2
XFILLER_235_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17388__A1 _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19453_ _18182_/B VGND VGND VPWR VPWR _19453_/Y sky130_fd_sc_hd__inv_2
X_16665_ _16664_/Y _16660_/X _16306_/X _16660_/X VGND VGND VPWR VPWR _16665_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _13861_/X _13875_/X _25197_/Q _13876_/X VGND VGND VPWR VPWR _13877_/X sky130_fd_sc_hd__o22a_4
XFILLER_222_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18404_ _16233_/Y _24179_/Q _16233_/Y _24179_/Q VGND VGND VPWR VPWR _18411_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15616_ _15616_/A VGND VGND VPWR VPWR _22651_/A sky130_fd_sc_hd__inv_2
X_12828_ _12828_/A VGND VGND VPWR VPWR _12828_/X sky130_fd_sc_hd__buf_2
X_19384_ _19381_/Y _19382_/X _19383_/X _19382_/X VGND VGND VPWR VPWR _19384_/X sky130_fd_sc_hd__a2bb2o_4
X_16596_ _24534_/Q VGND VGND VPWR VPWR _16596_/Y sky130_fd_sc_hd__inv_2
X_18335_ _18335_/A VGND VGND VPWR VPWR _20079_/B sky130_fd_sc_hd__buf_2
X_15547_ _15544_/A VGND VGND VPWR VPWR _15547_/X sky130_fd_sc_hd__buf_2
X_12759_ _12850_/A _23119_/A _12850_/A _23119_/A VGND VGND VPWR VPWR _12760_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18266_ _13828_/D _18262_/X _16090_/X _24231_/Q _18248_/A VGND VGND VPWR VPWR _24231_/D
+ sky130_fd_sc_hd__a32o_4
X_15478_ _15476_/Y _15472_/X _14427_/X _15477_/X VGND VGND VPWR VPWR _15478_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15083__A1_N _15082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17217_ _24618_/Q _17391_/A _24622_/Q _17358_/C VGND VGND VPWR VPWR _17220_/B sky130_fd_sc_hd__a2bb2o_4
X_14429_ _14425_/Y _14418_/X _14427_/X _14428_/X VGND VGND VPWR VPWR _14429_/X sky130_fd_sc_hd__a2bb2o_4
X_18197_ _18165_/A _19183_/A VGND VGND VPWR VPWR _18198_/C sky130_fd_sc_hd__or2_4
XFILLER_162_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17148_ _17127_/X _17144_/X _17148_/C VGND VGND VPWR VPWR _17148_/X sky130_fd_sc_hd__and3_4
X_17079_ _17079_/A VGND VGND VPWR VPWR _17080_/B sky130_fd_sc_hd__inv_2
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24129__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20090_ _13357_/B VGND VGND VPWR VPWR _20090_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24915__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16823__B1 _15738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22800_ _22535_/B VGND VGND VPWR VPWR _23072_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_20_0_HCLK clkbuf_7_10_0_HCLK/X VGND VGND VPWR VPWR _25543_/CLK sky130_fd_sc_hd__clkbuf_1
X_23780_ _23836_/CLK _23780_/D VGND VGND VPWR VPWR _17943_/B sky130_fd_sc_hd__dfxtp_4
X_20992_ _24129_/Q _24127_/Q VGND VGND VPWR VPWR _20992_/X sky130_fd_sc_hd__and2_4
XANTENNA__22947__A _22947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_83_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24812_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_226_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22731_ _16140_/Y _22444_/X _22730_/X _11811_/Y _22289_/X VGND VGND VPWR VPWR _22731_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25450_ _25454_/CLK _12475_/Y HRESETn VGND VGND VPWR VPWR _25450_/Q sky130_fd_sc_hd__dfrtp_4
X_22662_ _24630_/Q _22662_/B VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__or2_4
XFILLER_197_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20467__A _14550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24401_ _24952_/CLK _17095_/X HRESETn VGND VGND VPWR VPWR _24401_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22124__B2 _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21613_ _22226_/A VGND VGND VPWR VPWR _21644_/A sky130_fd_sc_hd__buf_2
X_25381_ _25380_/CLK _25381_/D HRESETn VGND VGND VPWR VPWR _25381_/Q sky130_fd_sc_hd__dfrtp_4
X_22593_ _21386_/B VGND VGND VPWR VPWR _22706_/B sky130_fd_sc_hd__buf_2
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_240_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24332_ _24334_/CLK _17444_/X HRESETn VGND VGND VPWR VPWR _24332_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21544_ _21544_/A _22897_/A VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__or2_4
XANTENNA__21883__B1 _24864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24263_ _24327_/CLK _24263_/D HRESETn VGND VGND VPWR VPWR _21066_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23085__C1 _23084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21475_ _18314_/X VGND VGND VPWR VPWR _21476_/A sky130_fd_sc_hd__buf_2
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23214_ _23137_/X _23212_/X _23139_/X _23213_/X VGND VGND VPWR VPWR _23215_/B sky130_fd_sc_hd__o22a_4
X_20426_ _20425_/Y _20423_/X _11847_/A _20423_/X VGND VGND VPWR VPWR _20426_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24194_ _24194_/CLK _24194_/D HRESETn VGND VGND VPWR VPWR _18490_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23145_ _20804_/Y _23006_/X _20943_/Y _22808_/X VGND VGND VPWR VPWR _23145_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13809__A _14412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20357_ _20356_/Y _20352_/X _20249_/X _20352_/X VGND VGND VPWR VPWR _23422_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23076_ _23076_/A _23183_/B VGND VGND VPWR VPWR _23076_/X sky130_fd_sc_hd__or2_4
X_20288_ _23448_/Q VGND VGND VPWR VPWR _21787_/B sky130_fd_sc_hd__inv_2
XFILLER_103_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22027_ _22027_/A VGND VGND VPWR VPWR _22028_/A sky130_fd_sc_hd__buf_2
XANTENNA__24656__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12570__A2_N _12568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16814__B1 HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13800_ _19595_/A _14264_/A VGND VGND VPWR VPWR _18268_/A sky130_fd_sc_hd__or2_4
XFILLER_229_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11992_ _11663_/B _11985_/X VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__and2_4
X_14780_ _14789_/A _14772_/C _14790_/B VGND VGND VPWR VPWR _14780_/X sky130_fd_sc_hd__o21a_4
XFILLER_217_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23978_ _23980_/CLK _23978_/D HRESETn VGND VGND VPWR VPWR _23978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13731_ _13695_/X _13729_/Y _13730_/X _13723_/X _11672_/A VGND VGND VPWR VPWR _25292_/D
+ sky130_fd_sc_hd__a32o_4
X_22929_ _21324_/X VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__buf_2
XFILLER_189_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16450_ HWDATA[2] VGND VGND VPWR VPWR _19091_/A sky130_fd_sc_hd__buf_2
XANTENNA__16886__A2_N _16877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13662_ _13660_/Y _13662_/B VGND VGND VPWR VPWR _13662_/X sky130_fd_sc_hd__and2_4
X_15401_ _15401_/A _15401_/B VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__or2_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12613_ _12613_/A VGND VGND VPWR VPWR _12710_/B sky130_fd_sc_hd__inv_2
X_13593_ _13593_/A VGND VGND VPWR VPWR _14569_/B sky130_fd_sc_hd__inv_2
X_16381_ _16381_/A VGND VGND VPWR VPWR _16382_/B sky130_fd_sc_hd__buf_2
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12603__B2 _24864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ _17984_/A _19470_/A VGND VGND VPWR VPWR _18120_/X sky130_fd_sc_hd__or2_4
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20677__A1 _14235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12544_ _25414_/Q VGND VGND VPWR VPWR _12725_/A sky130_fd_sc_hd__inv_2
X_15332_ _15318_/C _15329_/X VGND VGND VPWR VPWR _15332_/X sky130_fd_sc_hd__or2_4
XFILLER_129_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22592__A _22592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18051_ _18051_/A VGND VGND VPWR VPWR _18131_/A sky130_fd_sc_hd__buf_2
X_12475_ _12475_/A VGND VGND VPWR VPWR _12475_/Y sky130_fd_sc_hd__inv_2
X_15263_ _14895_/X _15260_/X VGND VGND VPWR VPWR _15264_/C sky130_fd_sc_hd__or2_4
XFILLER_185_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17002_ _17002_/A VGND VGND VPWR VPWR _17053_/C sky130_fd_sc_hd__inv_2
XFILLER_177_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14214_ _14214_/A VGND VGND VPWR VPWR _20525_/A sky130_fd_sc_hd__inv_2
X_15194_ _15193_/X VGND VGND VPWR VPWR _15195_/B sky130_fd_sc_hd__inv_2
XFILLER_126_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14145_ _14117_/X VGND VGND VPWR VPWR _14145_/X sky130_fd_sc_hd__buf_2
XFILLER_141_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12119__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14076_ _14058_/C _14074_/X _14066_/X _14008_/X _14075_/X VGND VGND VPWR VPWR _14076_/X
+ sky130_fd_sc_hd__a32o_4
X_18953_ _18951_/Y _18952_/X _16861_/X _18952_/X VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13027_ _13021_/A _13026_/X _13019_/A _13022_/Y VGND VGND VPWR VPWR _13027_/X sky130_fd_sc_hd__a211o_4
X_17904_ _17903_/Y _17913_/B _22003_/A _17901_/Y VGND VGND VPWR VPWR _17904_/X sky130_fd_sc_hd__o22a_4
X_18884_ _23957_/Q _20588_/B VGND VGND VPWR VPWR _18885_/B sky130_fd_sc_hd__or2_4
XANTENNA__24397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18310__A _21675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ _17832_/B VGND VGND VPWR VPWR _17836_/B sky130_fd_sc_hd__inv_2
XANTENNA__15653__B _11740_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17766_ _17766_/A _17766_/B _17824_/A _16950_/Y VGND VGND VPWR VPWR _17766_/X sky130_fd_sc_hd__or4_4
X_14978_ _14978_/A VGND VGND VPWR VPWR _14978_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19505_ _18289_/A _18288_/X _17723_/X VGND VGND VPWR VPWR _19505_/X sky130_fd_sc_hd__or3_4
XFILLER_207_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16717_ _16715_/Y _16716_/X _16537_/X _16716_/X VGND VGND VPWR VPWR _24489_/D sky130_fd_sc_hd__a2bb2o_4
X_13929_ _13929_/A VGND VGND VPWR VPWR _13951_/B sky130_fd_sc_hd__buf_2
X_17697_ _17696_/X VGND VGND VPWR VPWR _24300_/D sky130_fd_sc_hd__inv_2
X_19436_ _19166_/A _19436_/B _14665_/Y _13634_/X VGND VGND VPWR VPWR _19436_/X sky130_fd_sc_hd__or4_4
XFILLER_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16648_ _24516_/Q _16647_/X _16643_/X VGND VGND VPWR VPWR _24516_/D sky130_fd_sc_hd__o21a_4
XFILLER_222_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19367_ _19054_/A _19346_/B _19028_/C VGND VGND VPWR VPWR _19368_/A sky130_fd_sc_hd__or3_4
X_16579_ _16584_/A VGND VGND VPWR VPWR _16579_/X sky130_fd_sc_hd__buf_2
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22657__A2 _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18318_ _17743_/A VGND VGND VPWR VPWR _18325_/A sky130_fd_sc_hd__inv_2
XFILLER_194_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19298_ _21253_/B _19293_/X _18934_/X _19280_/Y VGND VGND VPWR VPWR _19298_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12517__B _13049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18249_ _18245_/X _18247_/X _16241_/A _22707_/A _18248_/X VGND VGND VPWR VPWR _24245_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21260_ _21260_/A _21257_/X _21260_/C VGND VGND VPWR VPWR _21260_/X sky130_fd_sc_hd__and3_4
X_20211_ _20211_/A VGND VGND VPWR VPWR _20211_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17297__B1 _17245_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21093__A1 _24786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21191_ _21182_/A VGND VGND VPWR VPWR _21211_/A sky130_fd_sc_hd__buf_2
X_20142_ _21629_/B _20141_/X _20119_/X _20141_/X VGND VGND VPWR VPWR _23503_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13858__B1 _13819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20073_ _20071_/Y _20072_/X _19807_/X _20072_/X VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__a2bb2o_4
X_24950_ _25103_/CLK _15506_/X HRESETn VGND VGND VPWR VPWR _11721_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18220__A _13639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23901_ _23885_/CLK _23901_/D VGND VGND VPWR VPWR _23901_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_246_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24881_ _24889_/CLK _24881_/D HRESETn VGND VGND VPWR VPWR _12535_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23832_ _23830_/CLK _19201_/X VGND VGND VPWR VPWR _19200_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_85_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14283__B1 _14248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22677__A _17257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23763_ _25077_/CLK _23763_/D VGND VGND VPWR VPWR _19394_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_72_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20975_ _12006_/B _13529_/A VGND VGND VPWR VPWR _24107_/D sky130_fd_sc_hd__and2_4
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25502_ _23615_/CLK _25502_/D HRESETn VGND VGND VPWR VPWR _11663_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_213_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22714_ _24433_/Q _22424_/B _15676_/A _22713_/X VGND VGND VPWR VPWR _22714_/X sky130_fd_sc_hd__a211o_4
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23694_ _23717_/CLK _19590_/X VGND VGND VPWR VPWR _23694_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16902__A1_N _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22645_ _22494_/X _22644_/X _21303_/A _24837_/Q _22569_/X VGND VGND VPWR VPWR _22645_/X
+ sky130_fd_sc_hd__a32o_4
X_25433_ _25433_/CLK _25433_/D HRESETn VGND VGND VPWR VPWR _25433_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15783__B1 _24860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25364_ _25358_/CLK _13044_/X HRESETn VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_139_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21856__B1 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22576_ _22562_/X _22574_/X _22144_/A _25535_/Q _22940_/A VGND VGND VPWR VPWR _22576_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_167_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21527_ _21512_/Y _21524_/Y _21526_/X VGND VGND VPWR VPWR _21527_/X sky130_fd_sc_hd__o21a_4
X_24315_ _24327_/CLK _17648_/X HRESETn VGND VGND VPWR VPWR _24315_/Q sky130_fd_sc_hd__dfrtp_4
X_25295_ _25292_/CLK _25295_/D HRESETn VGND VGND VPWR VPWR _11700_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ _12260_/A _12260_/B _12256_/X _12259_/X VGND VGND VPWR VPWR _12281_/B sky130_fd_sc_hd__or4_4
X_24246_ _24240_/CLK _24246_/D HRESETn VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21458_ _15792_/X VGND VGND VPWR VPWR _22447_/A sky130_fd_sc_hd__buf_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20409_ _20408_/X _20404_/X _11847_/A _23402_/Q _20406_/X VGND VGND VPWR VPWR _23402_/D
+ sky130_fd_sc_hd__a32o_4
X_12191_ _12191_/A VGND VGND VPWR VPWR _12191_/Y sky130_fd_sc_hd__inv_2
X_24177_ _23973_/CLK _24177_/D HRESETn VGND VGND VPWR VPWR _24177_/Q sky130_fd_sc_hd__dfrtp_4
X_21389_ _14688_/X _19853_/Y VGND VGND VPWR VPWR _21392_/B sky130_fd_sc_hd__or2_4
XANTENNA__24837__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23128_ _24711_/Q _22882_/X VGND VGND VPWR VPWR _23128_/X sky130_fd_sc_hd__or2_4
XFILLER_150_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15754__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15950_ HWDATA[28] VGND VGND VPWR VPWR _15950_/X sky130_fd_sc_hd__buf_2
X_23059_ _22788_/X _23057_/X _23058_/X _24744_/Q _22990_/X VGND VGND VPWR VPWR _23060_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19226__A _19091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14901_ _25019_/Q _14899_/Y _15196_/A _14914_/A VGND VGND VPWR VPWR _14901_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15881_ _12768_/Y _15877_/X _11766_/X _15880_/X VGND VGND VPWR VPWR _15881_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17620_ _17620_/A VGND VGND VPWR VPWR _17620_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13274__A _13420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14832_ _14832_/A _14837_/A VGND VGND VPWR VPWR _14832_/X sky130_fd_sc_hd__and2_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14274__B1 _13849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22587__A _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21491__A _22271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17551_ _24316_/Q VGND VGND VPWR VPWR _17579_/B sky130_fd_sc_hd__inv_2
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14763_ _21630_/A _14761_/X _14762_/Y VGND VGND VPWR VPWR _14763_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11975_ _25506_/Q _25505_/Q _11974_/X VGND VGND VPWR VPWR _11975_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19599__C _19550_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16502_ _24570_/Q VGND VGND VPWR VPWR _16502_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ _13702_/A _13702_/B VGND VGND VPWR VPWR _13714_/X sky130_fd_sc_hd__or2_4
XFILLER_17_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17482_ _18938_/B _17474_/X VGND VGND VPWR VPWR _17482_/Y sky130_fd_sc_hd__nor2_4
X_14694_ _14686_/X _14692_/B _14693_/Y VGND VGND VPWR VPWR _14695_/B sky130_fd_sc_hd__o21a_4
X_19221_ _19219_/Y _19217_/X _19220_/X _19217_/X VGND VGND VPWR VPWR _19221_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16433_ _16432_/Y _16428_/X _16248_/X _16428_/X VGND VGND VPWR VPWR _24597_/D sky130_fd_sc_hd__a2bb2o_4
X_13645_ _13644_/X VGND VGND VPWR VPWR _13645_/X sky130_fd_sc_hd__buf_2
XANTENNA__22639__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19152_ _19159_/A VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__buf_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16364_ _14400_/A VGND VGND VPWR VPWR _16364_/X sky130_fd_sc_hd__buf_2
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _25262_/Q _13575_/A _13574_/Y _13575_/Y VGND VGND VPWR VPWR _13587_/A sky130_fd_sc_hd__o22a_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _18199_/A _23833_/Q VGND VGND VPWR VPWR _18103_/X sky130_fd_sc_hd__or2_4
XFILLER_200_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15315_ _15307_/X _15314_/X VGND VGND VPWR VPWR _15315_/X sky130_fd_sc_hd__or2_4
XFILLER_157_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12527_ _12616_/A _24885_/Q _12616_/A _24885_/Q VGND VGND VPWR VPWR _12527_/X sky130_fd_sc_hd__a2bb2o_4
X_19083_ _19081_/Y _19077_/X _19012_/X _19082_/X VGND VGND VPWR VPWR _23874_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16295_ _16293_/Y _16291_/X _16294_/X _16291_/X VGND VGND VPWR VPWR _24647_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18034_ _17977_/A _23770_/Q VGND VGND VPWR VPWR _18037_/B sky130_fd_sc_hd__or2_4
X_15246_ _15245_/X VGND VGND VPWR VPWR _15246_/Y sky130_fd_sc_hd__inv_2
X_12458_ _12458_/A _12453_/X _12457_/X VGND VGND VPWR VPWR _25455_/D sky130_fd_sc_hd__and3_4
XFILLER_99_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12389_ _12382_/X _12384_/X _12389_/C _12388_/X VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__or4_4
X_15177_ _14897_/A _15176_/Y VGND VGND VPWR VPWR _15177_/X sky130_fd_sc_hd__or2_4
XFILLER_125_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12353__A _12353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24578__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14128_ _14121_/Y _14128_/B _14128_/C VGND VGND VPWR VPWR _14128_/X sky130_fd_sc_hd__and3_4
XFILLER_125_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19985_ _23556_/Q VGND VGND VPWR VPWR _22366_/B sky130_fd_sc_hd__inv_2
XANTENNA__24507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14059_ _14554_/A _14059_/B _14055_/Y _14058_/X VGND VGND VPWR VPWR _14059_/X sky130_fd_sc_hd__or4_4
X_18936_ _23924_/Q VGND VGND VPWR VPWR _18936_/Y sky130_fd_sc_hd__inv_2
X_18867_ _16519_/Y _18604_/X _24556_/Q _18685_/Y VGND VGND VPWR VPWR _18867_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18975__A _19091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17818_ _17762_/Y _17763_/Y _17562_/X _17761_/X VGND VGND VPWR VPWR _17818_/X sky130_fd_sc_hd__or4_4
XFILLER_239_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18798_ _18806_/A _18796_/X _18797_/X VGND VGND VPWR VPWR _24142_/D sky130_fd_sc_hd__and3_4
XFILLER_223_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17749_ _24293_/Q VGND VGND VPWR VPWR _17775_/C sky130_fd_sc_hd__inv_2
XANTENNA__16495__A _16495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20760_ _20739_/X _20759_/X _15611_/A _20744_/X VGND VGND VPWR VPWR _24029_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19419_ _19417_/Y _19415_/X _19418_/X _19415_/X VGND VGND VPWR VPWR _23755_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20691_ _20621_/B _20519_/X VGND VGND VPWR VPWR _24010_/D sky130_fd_sc_hd__and2_4
Xclkbuf_8_157_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24201_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22430_ _22430_/A _22430_/B VGND VGND VPWR VPWR _22430_/X sky130_fd_sc_hd__and2_4
XFILLER_149_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22361_ _22032_/A _19622_/Y VGND VGND VPWR VPWR _22362_/C sky130_fd_sc_hd__or2_4
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24100_ _24100_/CLK _20970_/X HRESETn VGND VGND VPWR VPWR RsTx_S0 sky130_fd_sc_hd__dfstp_4
XANTENNA__18215__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21312_ _24618_/Q _21312_/B VGND VGND VPWR VPWR _21312_/X sky130_fd_sc_hd__or2_4
XFILLER_248_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25080_ _25077_/CLK _25080_/D HRESETn VGND VGND VPWR VPWR _25080_/Q sky130_fd_sc_hd__dfrtp_4
X_22292_ _22289_/X _22291_/X _21308_/C _24727_/Q _21085_/X VGND VGND VPWR VPWR _22292_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22960__A _22836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24031_ _24495_/CLK _20770_/X HRESETn VGND VGND VPWR VPWR _20768_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21243_ _21267_/A _21243_/B VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__or2_4
XFILLER_190_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12263__A _25442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21576__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21174_ _16801_/Y _21592_/A _21332_/A _21173_/X VGND VGND VPWR VPWR _21174_/X sky130_fd_sc_hd__a211o_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20125_ _20124_/Y _20118_/X _19856_/X _20100_/Y VGND VGND VPWR VPWR _20125_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_22_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22566__A1 _22563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22566__B2 _22565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20056_ _20055_/Y _20051_/X _20034_/X _20038_/Y VGND VGND VPWR VPWR _23533_/D sky130_fd_sc_hd__a2bb2o_4
X_24933_ _24354_/CLK _24933_/D HRESETn VGND VGND VPWR VPWR _12077_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17442__B1 _16861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24864_ _24872_/CLK _15776_/X HRESETn VGND VGND VPWR VPWR _24864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23815_ _23454_/CLK _23815_/D VGND VGND VPWR VPWR _13381_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _24799_/CLK _24795_/D HRESETn VGND VGND VPWR VPWR _22139_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11759_/X VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_53_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20956_/A _20952_/A _20957_/X VGND VGND VPWR VPWR _20958_/Y sky130_fd_sc_hd__a21oi_4
X_23746_ _23669_/CLK _19445_/X VGND VGND VPWR VPWR _18044_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11691_/A VGND VGND VPWR VPWR _13690_/A sky130_fd_sc_hd__inv_2
XFILLER_199_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _13671_/A _13671_/B _20888_/Y VGND VGND VPWR VPWR _20889_/Y sky130_fd_sc_hd__a21oi_4
X_23677_ _24217_/CLK _19649_/X VGND VGND VPWR VPWR _19648_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21740__A2_N _16192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22854__B _22854_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13290_/X _13430_/B _13429_/X VGND VGND VPWR VPWR _13430_/X sky130_fd_sc_hd__and3_4
X_25416_ _25419_/CLK _12722_/X HRESETn VGND VGND VPWR VPWR _12622_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _16843_/A _22541_/X _22542_/X _22627_/X VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__a211o_4
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13286_/X _13361_/B VGND VGND VPWR VPWR _13361_/X sky130_fd_sc_hd__or2_4
X_22559_ _16522_/A _22440_/X _22545_/X VGND VGND VPWR VPWR _22559_/X sky130_fd_sc_hd__o21a_4
X_25347_ _25368_/CLK _13106_/X HRESETn VGND VGND VPWR VPWR _25347_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15100_ _25002_/Q _15098_/Y _25008_/Q _15099_/Y VGND VGND VPWR VPWR _15100_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23388__D HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12312_ _12311_/Y VGND VGND VPWR VPWR _12312_/X sky130_fd_sc_hd__buf_2
XFILLER_182_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13292_ _13468_/A _13292_/B VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__or2_4
X_16080_ _24723_/Q VGND VGND VPWR VPWR _16080_/Y sky130_fd_sc_hd__inv_2
X_25278_ _25276_/CLK _25278_/D HRESETn VGND VGND VPWR VPWR _25278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22870__A _22832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12243_ _25450_/Q VGND VGND VPWR VPWR _12296_/B sky130_fd_sc_hd__inv_2
X_15031_ _15005_/X _15011_/X _15021_/X _15031_/D VGND VGND VPWR VPWR _15031_/X sky130_fd_sc_hd__or4_4
X_24229_ _24230_/CLK _18272_/X HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24671__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12174_ _14359_/A VGND VGND VPWR VPWR _14334_/A sky130_fd_sc_hd__inv_2
XANTENNA__24600__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ _19768_/Y _19766_/X _19769_/X _19766_/X VGND VGND VPWR VPWR _19770_/X sky130_fd_sc_hd__a2bb2o_4
X_16982_ _24740_/Q _24397_/Q _16035_/Y _16981_/Y VGND VGND VPWR VPWR _16982_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14495__B1 _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18721_ _18739_/A _18719_/X _18720_/X VGND VGND VPWR VPWR _24160_/D sky130_fd_sc_hd__and3_4
XFILLER_107_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15933_ _19761_/A VGND VGND VPWR VPWR _15933_/X sky130_fd_sc_hd__buf_2
XFILLER_49_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18652_ _18645_/X _18649_/X _18650_/X _18651_/X VGND VGND VPWR VPWR _18652_/X sky130_fd_sc_hd__or4_4
XFILLER_67_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15864_ _15863_/X VGND VGND VPWR VPWR _15895_/A sky130_fd_sc_hd__buf_2
XANTENNA__22309__A1 _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17603_ _17663_/A _17594_/D VGND VGND VPWR VPWR _17616_/B sky130_fd_sc_hd__or2_4
XFILLER_236_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14815_ _14806_/Y _14815_/B _14815_/C VGND VGND VPWR VPWR _14816_/C sky130_fd_sc_hd__and3_4
X_18583_ _18556_/X _18570_/X _18582_/Y VGND VGND VPWR VPWR _24170_/D sky130_fd_sc_hd__and3_4
XANTENNA__15931__B _15934_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15795_ _15934_/B VGND VGND VPWR VPWR _15844_/A sky130_fd_sc_hd__inv_2
X_17534_ _17507_/X _17515_/X _17524_/X _17533_/X VGND VGND VPWR VPWR _17562_/A sky130_fd_sc_hd__or4_4
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ _14742_/Y _14745_/Y _14742_/A _14744_/X VGND VGND VPWR VPWR _14746_/X sky130_fd_sc_hd__o22a_4
X_11958_ _11955_/Y _11956_/X _11957_/X _11956_/X VGND VGND VPWR VPWR _11958_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17465_ _17463_/X _13306_/A _17464_/Y _13186_/Y VGND VGND VPWR VPWR _17465_/X sky130_fd_sc_hd__o22a_4
XFILLER_199_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15747__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14677_ _14668_/A _14676_/X _19028_/B _13610_/X VGND VGND VPWR VPWR _25078_/D sky130_fd_sc_hd__o22a_4
XFILLER_199_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11889_ _11889_/A VGND VGND VPWR VPWR _11889_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19204_ _19202_/Y _19203_/X _19091_/X _19203_/X VGND VGND VPWR VPWR _19204_/X sky130_fd_sc_hd__a2bb2o_4
X_16416_ _15105_/Y _16409_/X _16414_/X _16415_/X VGND VGND VPWR VPWR _24604_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13628_ _13628_/A _13628_/B VGND VGND VPWR VPWR _13628_/X sky130_fd_sc_hd__or2_4
X_17396_ _17396_/A VGND VGND VPWR VPWR _17396_/X sky130_fd_sc_hd__buf_2
XANTENNA__15762__A3 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19135_ _19133_/Y _19134_/X _19091_/X _19134_/X VGND VGND VPWR VPWR _19135_/X sky130_fd_sc_hd__a2bb2o_4
X_16347_ _16345_/Y _16346_/X _16252_/X _16346_/X VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__a2bb2o_4
X_13559_ _25266_/Q _14607_/A _13558_/Y _25092_/Q VGND VGND VPWR VPWR _13563_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24759__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12981__B1 _12875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19066_ _19065_/Y _19061_/X _18991_/X _19061_/X VGND VGND VPWR VPWR _23880_/D sky130_fd_sc_hd__a2bb2o_4
X_16278_ _16278_/A VGND VGND VPWR VPWR _16278_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16172__B1 _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18017_ _18097_/A VGND VGND VPWR VPWR _18063_/A sky130_fd_sc_hd__buf_2
X_15229_ _14935_/X _15228_/X _15183_/X VGND VGND VPWR VPWR _15229_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19968_ _22353_/B _19967_/X _19626_/X _19967_/X VGND VGND VPWR VPWR _23564_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14486__B1 _14420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22004__B _21991_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18919_ _23931_/Q VGND VGND VPWR VPWR _18919_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19899_ _23589_/Q VGND VGND VPWR VPWR _19899_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21930_ _21212_/A VGND VGND VPWR VPWR _21949_/A sky130_fd_sc_hd__buf_2
XANTENNA__25547__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21861_ _21861_/A VGND VGND VPWR VPWR _22176_/B sky130_fd_sc_hd__buf_2
XFILLER_103_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20812_ _20788_/X _20811_/X _15581_/A _20792_/X VGND VGND VPWR VPWR _20812_/X sky130_fd_sc_hd__a2bb2o_4
X_23600_ _23488_/CLK _23600_/D VGND VGND VPWR VPWR _23600_/Q sky130_fd_sc_hd__dfxtp_4
X_21792_ _21611_/X _21790_/X _21792_/C VGND VGND VPWR VPWR _21792_/X sky130_fd_sc_hd__and3_4
X_24580_ _24562_/CLK _16479_/X HRESETn VGND VGND VPWR VPWR _16478_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20743_ _20765_/A VGND VGND VPWR VPWR _20744_/A sky130_fd_sc_hd__buf_2
X_23531_ _23514_/CLK _20063_/X VGND VGND VPWR VPWR _23531_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _23669_/CLK _20252_/X VGND VGND VPWR VPWR _18178_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20674_ _17407_/A _17407_/B _20673_/Y _20622_/Y VGND VGND VPWR VPWR _20675_/C sky130_fd_sc_hd__a211o_4
XFILLER_184_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17768__B _17832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23276__A2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15753__A3 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22413_ _22413_/A _21069_/B VGND VGND VPWR VPWR _22413_/X sky130_fd_sc_hd__or2_4
X_25201_ _23998_/CLK _14246_/X HRESETn VGND VGND VPWR VPWR _25201_/Q sky130_fd_sc_hd__dfstp_4
X_23393_ _23913_/CLK _20426_/X VGND VGND VPWR VPWR _13229_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_164_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22344_ _21476_/A _22344_/B VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__or2_4
X_25132_ _25125_/CLK _14469_/X HRESETn VGND VGND VPWR VPWR _14467_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_148_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16163__B1 _16070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23028__A2 _21039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25063_ _24258_/CLK _14793_/X HRESETn VGND VGND VPWR VPWR _14785_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22275_ _22275_/A _19597_/X VGND VGND VPWR VPWR _22275_/X sky130_fd_sc_hd__and2_4
XANTENNA__15910__B1 _15629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24014_ _25106_/CLK _24014_/D HRESETn VGND VGND VPWR VPWR _24014_/Q sky130_fd_sc_hd__dfrtp_4
X_21226_ _21226_/A _21156_/X _21226_/C _21225_/X VGND VGND VPWR VPWR _21226_/X sky130_fd_sc_hd__and4_4
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21157_ _21157_/A _21375_/A VGND VGND VPWR VPWR _21157_/X sky130_fd_sc_hd__or2_4
XANTENNA__24011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20108_ _20108_/A VGND VGND VPWR VPWR _20108_/X sky130_fd_sc_hd__buf_2
XFILLER_219_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21088_ _22968_/B VGND VGND VPWR VPWR _23087_/B sky130_fd_sc_hd__buf_2
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12440__B _12247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12930_ _12927_/A _12926_/B _12929_/X VGND VGND VPWR VPWR _25390_/D sky130_fd_sc_hd__and3_4
X_20039_ _20038_/Y VGND VGND VPWR VPWR _20039_/X sky130_fd_sc_hd__buf_2
X_24916_ _24915_/CLK _15603_/X HRESETn VGND VGND VPWR VPWR _15601_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12856_/X _12860_/X VGND VGND VPWR VPWR _12895_/B sky130_fd_sc_hd__or2_4
X_24847_ _25425_/CLK _15817_/X HRESETn VGND VGND VPWR VPWR _24847_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14580_/Y _14595_/X _14598_/X _14599_/X _25098_/Q VGND VGND VPWR VPWR _14600_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13552__A _25265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ HWDATA[14] VGND VGND VPWR VPWR _16241_/A sky130_fd_sc_hd__buf_2
XPHY_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _23213_/A _15577_/X _11766_/X _15577_/X VGND VGND VPWR VPWR _24925_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17539__A1_N _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12790_/A _24819_/Q _12790_/Y _12791_/Y VGND VGND VPWR VPWR _12799_/B sky130_fd_sc_hd__o22a_4
X_24778_ _24803_/CLK _24778_/D HRESETn VGND VGND VPWR VPWR _24778_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15992__A3 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14531_ _25112_/Q _14520_/X _25111_/Q _14522_/X VGND VGND VPWR VPWR _14531_/X sky130_fd_sc_hd__o22a_4
XFILLER_199_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _15563_/A VGND VGND VPWR VPWR _21332_/A sky130_fd_sc_hd__inv_2
X_23729_ _23441_/CLK _19492_/X VGND VGND VPWR VPWR _19491_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16165__A1_N _16164_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15729__B1 _11763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17250_/A VGND VGND VPWR VPWR _17357_/A sky130_fd_sc_hd__inv_2
XFILLER_230_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14462_/A _14416_/X VGND VGND VPWR VPWR _14468_/A sky130_fd_sc_hd__nor2_4
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11672_/Y _24237_/Q _25301_/Q _22745_/A VGND VGND VPWR VPWR _11674_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14401__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_140_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23466_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16201_/A VGND VGND VPWR VPWR _16201_/Y sky130_fd_sc_hd__inv_2
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13413_/A _13413_/B VGND VGND VPWR VPWR _13413_/X sky130_fd_sc_hd__or2_4
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17181_ _17181_/A _17176_/X _17179_/X _17180_/X VGND VGND VPWR VPWR _17181_/X sky130_fd_sc_hd__or4_4
X_14393_ _14392_/X VGND VGND VPWR VPWR _14393_/X sky130_fd_sc_hd__buf_2
XFILLER_167_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14952__B2 _14954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24852__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16132_ _24703_/Q VGND VGND VPWR VPWR _16132_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11800__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13344_ _13207_/X _13343_/X _25335_/Q _13267_/X VGND VGND VPWR VPWR _25335_/D sky130_fd_sc_hd__o22a_4
XFILLER_194_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16063_ _24729_/Q VGND VGND VPWR VPWR _16063_/Y sky130_fd_sc_hd__inv_2
X_13275_ _13222_/X _13275_/B VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__or2_4
XANTENNA__15901__B1 _22641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15014_ _24480_/Q VGND VGND VPWR VPWR _15014_/Y sky130_fd_sc_hd__inv_2
X_12226_ _24782_/Q VGND VGND VPWR VPWR _12226_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22105__A _21879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12157_ _12157_/A VGND VGND VPWR VPWR _12157_/Y sky130_fd_sc_hd__inv_2
X_19822_ _19816_/A VGND VGND VPWR VPWR _19822_/X sky130_fd_sc_hd__buf_2
XFILLER_111_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16103__A _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12088_ _12083_/A VGND VGND VPWR VPWR _12088_/X sky130_fd_sc_hd__buf_2
X_16965_ _24718_/Q VGND VGND VPWR VPWR _16965_/Y sky130_fd_sc_hd__inv_2
X_19753_ _11861_/A VGND VGND VPWR VPWR _19753_/X sky130_fd_sc_hd__buf_2
X_15916_ _12797_/Y _15912_/X _15486_/X _15912_/X VGND VGND VPWR VPWR _24792_/D sky130_fd_sc_hd__a2bb2o_4
X_18704_ _18733_/C _18711_/A VGND VGND VPWR VPWR _18717_/B sky130_fd_sc_hd__or2_4
X_19684_ _13325_/B VGND VGND VPWR VPWR _19684_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19414__A _19413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16896_ _20146_/A VGND VGND VPWR VPWR _16896_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21753__A2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18635_ _24160_/Q VGND VGND VPWR VPWR _18720_/A sky130_fd_sc_hd__inv_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15847_ _12343_/Y _15842_/X _15486_/X _15842_/X VGND VGND VPWR VPWR _15847_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18566_ _18595_/A _18425_/Y _18433_/Y _18565_/X VGND VGND VPWR VPWR _18566_/X sky130_fd_sc_hd__or4_4
X_15778_ _15758_/X _15774_/X _15777_/X _24863_/Q _15719_/X VGND VGND VPWR VPWR _15778_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_206_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22775__A _22774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17517_ _25544_/Q _24315_/Q _11792_/Y _17516_/Y VGND VGND VPWR VPWR _17517_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14729_ _14729_/A VGND VGND VPWR VPWR _14729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17869__A _17861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18497_ _18488_/A _18487_/X VGND VGND VPWR VPWR _18510_/B sky130_fd_sc_hd__or2_4
XFILLER_32_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17448_ _17448_/A _17448_/B _17448_/C VGND VGND VPWR VPWR _17448_/X sky130_fd_sc_hd__or3_4
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15735__A3 _15734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22466__B1 _15108_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17379_ _17363_/A _17375_/X _17378_/Y VGND VGND VPWR VPWR _17379_/X sky130_fd_sc_hd__and3_4
XFILLER_229_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24593__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19118_ _13189_/B VGND VGND VPWR VPWR _19118_/Y sky130_fd_sc_hd__inv_2
X_20390_ _20390_/A VGND VGND VPWR VPWR _22045_/B sky130_fd_sc_hd__inv_2
XFILLER_145_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19049_ _19046_/Y _19044_/X _19048_/X _19044_/X VGND VGND VPWR VPWR _19049_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22769__A1 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22060_ _22060_/A _19610_/X VGND VGND VPWR VPWR _22060_/X sky130_fd_sc_hd__and2_4
XFILLER_160_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ _21010_/A _24343_/Q _24344_/Q _21010_/X VGND VGND VPWR VPWR _23984_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14459__B1 _14248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19398__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16948__A _24291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22962_ _12269_/Y _23280_/A _22961_/X VGND VGND VPWR VPWR _22962_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24701_ _24756_/CLK _16139_/X HRESETn VGND VGND VPWR VPWR _22763_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21913_ _14709_/X _21902_/X _21912_/X VGND VGND VPWR VPWR _21913_/X sky130_fd_sc_hd__or3_4
XFILLER_243_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22893_ _23072_/A _22893_/B VGND VGND VPWR VPWR _22893_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14468__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24632_ _24629_/CLK _24632_/D HRESETn VGND VGND VPWR VPWR _24632_/Q sky130_fd_sc_hd__dfrtp_4
X_21844_ _21040_/Y VGND VGND VPWR VPWR _21844_/X sky130_fd_sc_hd__buf_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21630_/A _21773_/X _21775_/C VGND VGND VPWR VPWR _21775_/X sky130_fd_sc_hd__and3_4
X_24563_ _24562_/CLK _16521_/X HRESETn VGND VGND VPWR VPWR _16519_/A sky130_fd_sc_hd__dfrtp_4
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _20725_/X VGND VGND VPWR VPWR _20731_/B sky130_fd_sc_hd__inv_2
X_23514_ _23514_/CLK _20110_/X VGND VGND VPWR VPWR _20107_/A sky130_fd_sc_hd__dfxtp_4
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24494_ _24493_/CLK _16705_/X HRESETn VGND VGND VPWR VPWR _24494_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20180__B2 _20177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_213_0_HCLK clkbuf_7_106_0_HCLK/X VGND VGND VPWR VPWR _25023_/CLK sky130_fd_sc_hd__clkbuf_1
X_20657_ _17404_/B _20656_/Y _20669_/C VGND VGND VPWR VPWR _20657_/X sky130_fd_sc_hd__and3_4
X_23445_ _23445_/CLK _20296_/X VGND VGND VPWR VPWR _23445_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23376_ _21002_/X VGND VGND VPWR VPWR IRQ[20] sky130_fd_sc_hd__buf_2
X_20588_ _23957_/Q _20588_/B VGND VGND VPWR VPWR _20588_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25115_ _23970_/CLK _25115_/D HRESETn VGND VGND VPWR VPWR _14510_/B sky130_fd_sc_hd__dfrtp_4
X_22327_ _22320_/Y _22322_/Y _22323_/X _22327_/D VGND VGND VPWR VPWR _22327_/X sky130_fd_sc_hd__or4_4
XFILLER_191_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ _13059_/X VGND VGND VPWR VPWR _25360_/D sky130_fd_sc_hd__inv_2
X_22258_ _18301_/A _22254_/X _22257_/X VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__or3_4
X_25046_ _24000_/CLK _25046_/D HRESETn VGND VGND VPWR VPWR _14889_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12011_ _12009_/A _12010_/A _12009_/Y _12010_/Y VGND VGND VPWR VPWR _12011_/X sky130_fd_sc_hd__o22a_4
X_21209_ _21209_/A _21209_/B _21208_/X VGND VGND VPWR VPWR _21209_/X sky130_fd_sc_hd__and3_4
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22189_ _22188_/X VGND VGND VPWR VPWR _22189_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23185__A1 _16482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16750_ _16750_/A VGND VGND VPWR VPWR _16750_/Y sky130_fd_sc_hd__inv_2
X_13962_ _13944_/A _15435_/B _13962_/C VGND VGND VPWR VPWR _13962_/X sky130_fd_sc_hd__or3_4
XFILLER_219_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15701_ _15701_/A _15701_/B VGND VGND VPWR VPWR _18029_/A sky130_fd_sc_hd__or2_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _12859_/X _12921_/D VGND VGND VPWR VPWR _12913_/X sky130_fd_sc_hd__or2_4
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16681_ _16679_/Y _16680_/X _16412_/X _16680_/X VGND VGND VPWR VPWR _24504_/D sky130_fd_sc_hd__a2bb2o_4
X_13893_ _23979_/Q VGND VGND VPWR VPWR _13893_/X sky130_fd_sc_hd__buf_2
XFILLER_206_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18420_ _18420_/A _18415_/X _18420_/C _18419_/X VGND VGND VPWR VPWR _18420_/X sky130_fd_sc_hd__or4_4
XFILLER_207_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13282__A _13282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15632_ _14423_/A VGND VGND VPWR VPWR _15632_/X sky130_fd_sc_hd__buf_2
X_12844_ _12838_/X _12840_/X _12844_/C _12843_/X VGND VGND VPWR VPWR _12845_/D sky130_fd_sc_hd__or4_4
X_18351_ _13198_/A _18349_/B VGND VGND VPWR VPWR _18351_/X sky130_fd_sc_hd__and2_4
X_15563_ _15563_/A VGND VGND VPWR VPWR _21172_/B sky130_fd_sc_hd__buf_2
XANTENNA__22696__B1 _21229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12775_ _12773_/A _22875_/A _12773_/Y _12774_/Y VGND VGND VPWR VPWR _12786_/A sky130_fd_sc_hd__o22a_4
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17248_/B _17301_/X VGND VGND VPWR VPWR _17305_/B sky130_fd_sc_hd__or2_4
XANTENNA__19561__B1 _19560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14514_ _14510_/C VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__buf_2
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _12061_/A VGND VGND VPWR VPWR _11727_/A sky130_fd_sc_hd__inv_2
X_18282_ _19527_/C VGND VGND VPWR VPWR _18282_/X sky130_fd_sc_hd__buf_2
XFILLER_202_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ HTRANS[1] VGND VGND VPWR VPWR _15494_/Y sky130_fd_sc_hd__inv_2
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _17226_/X _17233_/B _17233_/C _17232_/X VGND VGND VPWR VPWR _17233_/X sky130_fd_sc_hd__or4_4
X_14445_ _15471_/A _14388_/B VGND VGND VPWR VPWR _14446_/A sky130_fd_sc_hd__nor2_4
XFILLER_175_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22448__B1 _12327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11657_/A VGND VGND VPWR VPWR _11658_/A sky130_fd_sc_hd__inv_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22999__B2 _22924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _17137_/B _17163_/X VGND VGND VPWR VPWR _17166_/B sky130_fd_sc_hd__or2_4
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14364_/A _14375_/X _12092_/A _14369_/X VGND VGND VPWR VPWR _25162_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22463__A3 _16468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16115_ _24710_/Q VGND VGND VPWR VPWR _16115_/Y sky130_fd_sc_hd__inv_2
X_13327_ _13242_/X _13325_/X _13326_/X VGND VGND VPWR VPWR _13327_/X sky130_fd_sc_hd__and3_4
X_17095_ _17095_/A _17088_/B _17094_/X VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__and3_4
XFILLER_142_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16046_ _24736_/Q VGND VGND VPWR VPWR _16046_/Y sky130_fd_sc_hd__inv_2
X_13258_ _13257_/X _13258_/B VGND VGND VPWR VPWR _13258_/X sky130_fd_sc_hd__or2_4
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12209_ _22871_/A VGND VGND VPWR VPWR _12209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13457__A _13356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _13192_/A _13189_/B VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__or2_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19805_ _19805_/A VGND VGND VPWR VPWR _21621_/B sky130_fd_sc_hd__inv_2
XANTENNA__15102__B2 _24585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17997_ _18102_/A VGND VGND VPWR VPWR _18191_/A sky130_fd_sc_hd__buf_2
XFILLER_85_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15672__A _21170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16948_ _24291_/Q VGND VGND VPWR VPWR _16957_/A sky130_fd_sc_hd__inv_2
X_19736_ _13432_/B VGND VGND VPWR VPWR _19736_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_211_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16879_ _24415_/Q VGND VGND VPWR VPWR _19800_/A sky130_fd_sc_hd__buf_2
X_19667_ _19652_/Y VGND VGND VPWR VPWR _19667_/X sky130_fd_sc_hd__buf_2
XFILLER_237_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _18617_/Y VGND VGND VPWR VPWR _18756_/A sky130_fd_sc_hd__buf_2
XFILLER_52_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19598_ _19597_/X VGND VGND VPWR VPWR _19599_/D sky130_fd_sc_hd__buf_2
XFILLER_241_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15956__A3 HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17599__A _17691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18549_ _18543_/A _18543_/B VGND VGND VPWR VPWR _18549_/Y sky130_fd_sc_hd__nand2_4
XFILLER_178_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24774__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21560_ _21560_/A _22129_/B VGND VGND VPWR VPWR _21563_/B sky130_fd_sc_hd__nand2_4
XANTENNA__16366__B1 _16364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15169__B2 _24588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24703__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20511_ _20511_/A _20620_/A _20511_/C VGND VGND VPWR VPWR _20511_/X sky130_fd_sc_hd__and3_4
XFILLER_21_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21491_ _22271_/A VGND VGND VPWR VPWR _21688_/A sky130_fd_sc_hd__buf_2
X_23230_ _23321_/A _23229_/X VGND VGND VPWR VPWR _23230_/X sky130_fd_sc_hd__and2_4
XFILLER_193_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20442_ _20442_/A VGND VGND VPWR VPWR _20443_/B sky130_fd_sc_hd__inv_2
XFILLER_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23161_ _23117_/A _23160_/X VGND VGND VPWR VPWR _23161_/X sky130_fd_sc_hd__and2_4
XANTENNA__21662__A1 _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20373_ _20372_/Y _20370_/X _19636_/A _20370_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_43_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23516_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22112_ _20470_/A _22176_/B VGND VGND VPWR VPWR _22119_/A sky130_fd_sc_hd__nor2_4
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23092_ _24745_/Q _21039_/X _21068_/X _23091_/X VGND VGND VPWR VPWR _23093_/C sky130_fd_sc_hd__a211o_4
X_22043_ _22036_/A _22041_/X _22043_/C VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__and3_4
XFILLER_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23994_ _23998_/CLK _20659_/Y HRESETn VGND VGND VPWR VPWR _23994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_228_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22945_ _22945_/A VGND VGND VPWR VPWR _23189_/B sky130_fd_sc_hd__buf_2
XFILLER_216_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14629__C _14679_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22876_ _22488_/X _22875_/X _21434_/X _24878_/Q _22784_/X VGND VGND VPWR VPWR _22877_/B
+ sky130_fd_sc_hd__a32o_4
X_24615_ _24613_/CLK _24615_/D HRESETn VGND VGND VPWR VPWR _16387_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_231_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21827_ _21808_/A _21825_/X _21826_/X VGND VGND VPWR VPWR _21827_/X sky130_fd_sc_hd__and3_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _25408_/Q VGND VGND VPWR VPWR _12742_/A sky130_fd_sc_hd__inv_2
X_24546_ _24562_/CLK _24546_/D HRESETn VGND VGND VPWR VPWR _16566_/A sky130_fd_sc_hd__dfrtp_4
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16357__B1 _16066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12091__B1 _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23023__B _22954_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21758_ _21606_/A _21756_/X _21123_/A _21757_/X VGND VGND VPWR VPWR _21758_/X sky130_fd_sc_hd__o22a_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14460__A1_N _14191_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _20708_/Y _13132_/X _13134_/X VGND VGND VPWR VPWR _20709_/X sky130_fd_sc_hd__o21a_4
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12228_/A _12491_/B VGND VGND VPWR VPWR _12491_/X sky130_fd_sc_hd__or2_4
X_24477_ _24473_/CLK _16749_/X HRESETn VGND VGND VPWR VPWR _24477_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21689_ _22029_/A _21689_/B _21689_/C VGND VGND VPWR VPWR _21689_/X sky130_fd_sc_hd__and3_4
XFILLER_184_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _14230_/A VGND VGND VPWR VPWR _14232_/A sky130_fd_sc_hd__buf_2
XFILLER_138_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428_ _24217_/CLK _20341_/X VGND VGND VPWR VPWR _20340_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16109__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21759__A _21604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22445__A3 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14161_ _14153_/X _14160_/Y _14110_/A _14153_/X VGND VGND VPWR VPWR _25223_/D sky130_fd_sc_hd__a2bb2o_4
X_23359_ _24229_/Q _21997_/X _23357_/X _23358_/Y VGND VGND VPWR VPWR _23360_/B sky130_fd_sc_hd__a211o_4
XFILLER_165_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13112_ _13107_/B _13111_/X _13121_/C VGND VGND VPWR VPWR _25345_/D sky130_fd_sc_hd__and3_4
X_14092_ _14027_/B _14090_/X _14087_/X _14027_/A _14085_/X VGND VGND VPWR VPWR _25238_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13277__A _13315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13043_ _12329_/Y _13039_/B VGND VGND VPWR VPWR _13043_/Y sky130_fd_sc_hd__nand2_4
X_17920_ _17919_/Y _17915_/Y _22005_/A _17915_/A VGND VGND VPWR VPWR _24259_/D sky130_fd_sc_hd__o22a_4
X_25029_ _25030_/CLK _25029_/D HRESETn VGND VGND VPWR VPWR _25029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17851_ _17762_/Y _17849_/A VGND VGND VPWR VPWR _17851_/X sky130_fd_sc_hd__or2_4
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16588__A _24537_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16802_ _16801_/Y _16738_/X _16729_/X _16738_/X VGND VGND VPWR VPWR _16802_/X sky130_fd_sc_hd__a2bb2o_4
X_17782_ _16925_/Y _16957_/X _17781_/X VGND VGND VPWR VPWR _17782_/X sky130_fd_sc_hd__or3_4
X_14994_ _14994_/A _14994_/B VGND VGND VPWR VPWR _15067_/A sky130_fd_sc_hd__or2_4
XFILLER_226_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21169__B1 _21332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _16733_/A VGND VGND VPWR VPWR _22592_/A sky130_fd_sc_hd__buf_2
X_19521_ _21665_/B _19520_/X _11961_/X _19520_/X VGND VGND VPWR VPWR _23719_/D sky130_fd_sc_hd__a2bb2o_4
X_13945_ _13945_/A VGND VGND VPWR VPWR _14257_/D sky130_fd_sc_hd__inv_2
XFILLER_47_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14413__A1_N _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19452_ _19450_/Y _19451_/X _19383_/X _19451_/X VGND VGND VPWR VPWR _23743_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16664_ _16664_/A VGND VGND VPWR VPWR _16664_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13876_ _13876_/A VGND VGND VPWR VPWR _13876_/X sky130_fd_sc_hd__buf_2
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15615_ _15613_/Y _15609_/X _11818_/X _15614_/X VGND VGND VPWR VPWR _24911_/D sky130_fd_sc_hd__a2bb2o_4
X_18403_ _18398_/X _18399_/X _18401_/X _18402_/X VGND VGND VPWR VPWR _18403_/X sky130_fd_sc_hd__or4_4
XFILLER_62_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12827_ _25377_/Q VGND VGND VPWR VPWR _12828_/A sky130_fd_sc_hd__inv_2
X_19383_ _11865_/X VGND VGND VPWR VPWR _19383_/X sky130_fd_sc_hd__buf_2
XFILLER_50_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16595_ _16594_/Y _16592_/X _16238_/X _16592_/X VGND VGND VPWR VPWR _24535_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18334_ _17463_/X VGND VGND VPWR VPWR _18334_/X sky130_fd_sc_hd__buf_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17212__A _17212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15546_ _12107_/X _15544_/X HADDR[3] _15544_/X VGND VGND VPWR VPWR _24933_/D sky130_fd_sc_hd__a2bb2o_4
X_12758_ _12899_/A VGND VGND VPWR VPWR _12850_/A sky130_fd_sc_hd__inv_2
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20144__B2 _20141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A _11684_/X _11709_/C _11708_/X VGND VGND VPWR VPWR _11889_/A sky130_fd_sc_hd__or4_4
X_18265_ _11692_/Y _18243_/A _16726_/X _18243_/A VGND VGND VPWR VPWR _24232_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21892__A1 _25442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15477_ _15472_/A VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__buf_2
XANTENNA__24114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12689_ _12619_/B _12689_/B VGND VGND VPWR VPWR _12689_/X sky130_fd_sc_hd__or2_4
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _24351_/Q VGND VGND VPWR VPWR _17358_/C sky130_fd_sc_hd__inv_2
X_14428_ _14428_/A VGND VGND VPWR VPWR _14428_/X sky130_fd_sc_hd__buf_2
X_18196_ _18164_/A _19161_/A VGND VGND VPWR VPWR _18198_/B sky130_fd_sc_hd__or2_4
XANTENNA__23094__B1 _17753_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17866__B _17861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12385__B2 _24829_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17147_ _17050_/D _17143_/X VGND VGND VPWR VPWR _17148_/C sky130_fd_sc_hd__nand2_4
X_14359_ _14359_/A _14359_/B _14358_/X VGND VGND VPWR VPWR _14359_/X sky130_fd_sc_hd__and3_4
XANTENNA__19139__A _19139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_2_0_HCLK clkbuf_7_1_0_HCLK/X VGND VGND VPWR VPWR _23555_/CLK sky130_fd_sc_hd__clkbuf_1
X_17078_ _17078_/A VGND VGND VPWR VPWR _24406_/D sky130_fd_sc_hd__inv_2
XFILLER_226_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16029_ _16028_/Y _16024_/X _15960_/X _16024_/X VGND VGND VPWR VPWR _16029_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13187__A _13186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19719_ _19719_/A VGND VGND VPWR VPWR _19719_/Y sky130_fd_sc_hd__inv_2
X_20991_ _24126_/Q _24124_/Q _24125_/Q _20990_/X VGND VGND VPWR VPWR _20991_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22730_ _22284_/X VGND VGND VPWR VPWR _22730_/X sky130_fd_sc_hd__buf_2
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16587__B1 _16417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23124__A _22721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22661_ _22629_/X _22636_/Y _22640_/X _22660_/Y VGND VGND VPWR VPWR HRDATA[12] sky130_fd_sc_hd__or4_4
XFILLER_41_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18328__A1 _21834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22124__A2 _15792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24400_ _24952_/CLK _24400_/D HRESETn VGND VGND VPWR VPWR _17018_/A sky130_fd_sc_hd__dfrtp_4
X_21612_ _21263_/A VGND VGND VPWR VPWR _22226_/A sky130_fd_sc_hd__buf_2
XANTENNA__15648__A2_N _15584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25380_ _25380_/CLK _25380_/D HRESETn VGND VGND VPWR VPWR _25380_/Q sky130_fd_sc_hd__dfrtp_4
X_22592_ _22592_/A _22592_/B _22591_/X VGND VGND VPWR VPWR _22592_/X sky130_fd_sc_hd__and3_4
XFILLER_187_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20135__B2 _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24331_ _24334_/CLK _24331_/D HRESETn VGND VGND VPWR VPWR _17445_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21883__A1 _24794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21543_ _21543_/A VGND VGND VPWR VPWR _22897_/A sky130_fd_sc_hd__buf_2
XFILLER_178_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21883__B2 _21085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22682__B _21882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21474_ _21474_/A _21474_/B VGND VGND VPWR VPWR _21478_/B sky130_fd_sc_hd__or2_4
X_24262_ _23597_/CLK _24262_/D HRESETn VGND VGND VPWR VPWR _24262_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20425_ _13229_/B VGND VGND VPWR VPWR _20425_/Y sky130_fd_sc_hd__inv_2
X_23213_ _23213_/A _22890_/B VGND VGND VPWR VPWR _23213_/X sky130_fd_sc_hd__and2_4
XANTENNA__15577__A _15584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12376__B2 _12375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24193_ _24194_/CLK _18496_/Y HRESETn VGND VGND VPWR VPWR _24193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21298__B _21307_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20356_ _23422_/Q VGND VGND VPWR VPWR _20356_/Y sky130_fd_sc_hd__inv_2
X_23144_ _23144_/A VGND VGND VPWR VPWR _23249_/A sky130_fd_sc_hd__buf_2
XANTENNA__16511__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23075_ _22738_/A VGND VGND VPWR VPWR _23183_/B sky130_fd_sc_hd__buf_2
X_20287_ _21921_/B _20284_/X _19800_/A _20284_/X VGND VGND VPWR VPWR _23449_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22026_ _22034_/A _22026_/B VGND VGND VPWR VPWR _22029_/B sky130_fd_sc_hd__or2_4
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18264__B1 _16861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16201__A _16201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22899__B1 _22815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11991_ _11663_/C _11990_/X _11988_/X VGND VGND VPWR VPWR _11991_/X sky130_fd_sc_hd__o21a_4
X_23977_ _24334_/CLK _23977_/D HRESETn VGND VGND VPWR VPWR _20548_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__24696__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _13688_/Y VGND VGND VPWR VPWR _13730_/X sky130_fd_sc_hd__buf_2
XFILLER_216_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22928_ _17263_/C _22926_/X _25392_/Q _22927_/X VGND VGND VPWR VPWR _22928_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24625__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13661_ _24048_/Q _24047_/Q VGND VGND VPWR VPWR _13662_/B sky130_fd_sc_hd__nor2_4
X_22859_ _12237_/Y _22286_/X _16468_/A _12350_/Y _22858_/X VGND VGND VPWR VPWR _22859_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14656__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15400_ _15415_/A _15399_/X VGND VGND VPWR VPWR _15401_/B sky130_fd_sc_hd__or2_4
XFILLER_231_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12612_ _12730_/A VGND VGND VPWR VPWR _12636_/A sky130_fd_sc_hd__buf_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17032__A _24650_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16380_ _14199_/A _22459_/A VGND VGND VPWR VPWR _16381_/A sky130_fd_sc_hd__or2_4
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13592_ _13589_/Y _25098_/Q _25264_/Q _14613_/A VGND VGND VPWR VPWR _13596_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22666__A3 _22148_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15331_ _25010_/Q _15331_/B VGND VGND VPWR VPWR _15331_/X sky130_fd_sc_hd__or2_4
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12543_ _12541_/A _24879_/Q _12618_/A _12542_/Y VGND VGND VPWR VPWR _12543_/X sky130_fd_sc_hd__o22a_4
X_24529_ _24528_/CLK _16611_/X HRESETn VGND VGND VPWR VPWR _24529_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18050_ _17954_/A _18042_/X _18049_/X VGND VGND VPWR VPWR _18050_/X sky130_fd_sc_hd__and3_4
X_15262_ _25024_/Q _15261_/Y VGND VGND VPWR VPWR _15262_/X sky130_fd_sc_hd__or2_4
X_12474_ _12439_/B _12468_/X _12421_/A _12470_/Y VGND VGND VPWR VPWR _12475_/A sky130_fd_sc_hd__a211o_4
XFILLER_145_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17001_ _24738_/Q _17118_/A _16072_/Y _17159_/A VGND VGND VPWR VPWR _17001_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14213_ _20518_/A _14208_/X _13846_/X _14210_/X VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__a2bb2o_4
X_15193_ _15193_/A _15294_/A VGND VGND VPWR VPWR _15193_/X sky130_fd_sc_hd__or2_4
XANTENNA__25484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14144_ _14112_/A _14112_/B _14112_/A _14112_/B VGND VGND VPWR VPWR _14144_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_152_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14075_ _14069_/B VGND VGND VPWR VPWR _14075_/X sky130_fd_sc_hd__buf_2
X_18952_ _18952_/A VGND VGND VPWR VPWR _18952_/X sky130_fd_sc_hd__buf_2
XFILLER_113_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13026_ _13026_/A _13008_/X _13026_/C _13026_/D VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__or4_4
X_17903_ _22003_/A VGND VGND VPWR VPWR _17903_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22051__A1 _22274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15934__B _15934_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18883_ _20584_/A _18883_/B VGND VGND VPWR VPWR _20588_/B sky130_fd_sc_hd__or2_4
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17834_ _17852_/A _17834_/B _17833_/Y VGND VGND VPWR VPWR _24281_/D sky130_fd_sc_hd__and3_4
XFILLER_239_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15653__C _11740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18653__A1_N _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21952__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23000__B1 _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14977_ _15258_/A _24423_/Q _15002_/A _14976_/Y VGND VGND VPWR VPWR _14983_/B sky130_fd_sc_hd__a2bb2o_4
X_17765_ _24277_/Q VGND VGND VPWR VPWR _17766_/B sky130_fd_sc_hd__inv_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19504_ _18290_/A VGND VGND VPWR VPWR _19965_/A sky130_fd_sc_hd__buf_2
XANTENNA__15950__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13928_ _13928_/A VGND VGND VPWR VPWR _13951_/A sky130_fd_sc_hd__buf_2
X_16716_ _16709_/A VGND VGND VPWR VPWR _16716_/X sky130_fd_sc_hd__buf_2
X_17696_ _17588_/B _17672_/X _17693_/Y _17611_/X VGND VGND VPWR VPWR _17696_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16647_ _16182_/B _16633_/X VGND VGND VPWR VPWR _16647_/X sky130_fd_sc_hd__and2_4
X_19435_ _17963_/B VGND VGND VPWR VPWR _19435_/Y sky130_fd_sc_hd__inv_2
X_13859_ _24008_/Q VGND VGND VPWR VPWR _13872_/A sky130_fd_sc_hd__inv_2
XFILLER_222_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18668__A1_N _16625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18038__A _18006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16578_ _16578_/A VGND VGND VPWR VPWR _16578_/Y sky130_fd_sc_hd__inv_2
X_19366_ _17955_/B VGND VGND VPWR VPWR _19366_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15529_ _15528_/Y _15526_/X HADDR[11] _15526_/X VGND VGND VPWR VPWR _24941_/D sky130_fd_sc_hd__a2bb2o_4
X_18317_ _21676_/A _18297_/X _18310_/X VGND VGND VPWR VPWR _24217_/D sky130_fd_sc_hd__a21oi_4
XFILLER_175_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19297_ _19297_/A VGND VGND VPWR VPWR _21253_/B sky130_fd_sc_hd__inv_2
XFILLER_187_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ _18248_/A VGND VGND VPWR VPWR _18248_/X sky130_fd_sc_hd__buf_2
XFILLER_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23067__B1 _12817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16741__B1 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18179_ _17991_/X _18177_/X _18178_/X VGND VGND VPWR VPWR _18180_/C sky130_fd_sc_hd__and3_4
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20210_ _20209_/Y _20205_/X _20146_/X _20193_/A VGND VGND VPWR VPWR _23477_/D sky130_fd_sc_hd__a2bb2o_4
X_21190_ _21207_/A _21190_/B VGND VGND VPWR VPWR _21190_/X sky130_fd_sc_hd__or2_4
XFILLER_143_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20141_ _20129_/A VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__buf_2
XFILLER_144_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_117_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _25419_/CLK sky130_fd_sc_hd__clkbuf_1
X_20072_ _20059_/Y VGND VGND VPWR VPWR _20072_/X sky130_fd_sc_hd__buf_2
XFILLER_98_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23900_ _23885_/CLK _23900_/D VGND VGND VPWR VPWR _19001_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_218_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24880_ _24889_/CLK _15743_/X HRESETn VGND VGND VPWR VPWR _12593_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18261__A3 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23831_ _24100_/CLK _19204_/X VGND VGND VPWR VPWR _23831_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15860__A _21173_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22677__B _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23762_ _25077_/CLK _23762_/D VGND VGND VPWR VPWR _23762_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20974_ _12019_/A _13529_/A VGND VGND VPWR VPWR _24106_/D sky130_fd_sc_hd__and2_4
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25501_ _23615_/CLK _25501_/D HRESETn VGND VGND VPWR VPWR _11663_/B sky130_fd_sc_hd__dfrtp_4
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22713_ _22713_/A _21855_/B _21752_/B VGND VGND VPWR VPWR _22713_/X sky130_fd_sc_hd__and3_4
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23693_ _23717_/CLK _19592_/X VGND VGND VPWR VPWR _19591_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_213_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25432_ _25433_/CLK _25432_/D HRESETn VGND VGND VPWR VPWR _25432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22644_ _22644_/A _22789_/B VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__or2_4
XFILLER_201_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13794__B1 _13481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25363_ _25365_/CLK _13047_/X HRESETn VGND VGND VPWR VPWR _12363_/A sky130_fd_sc_hd__dfrtp_4
X_22575_ _22575_/A VGND VGND VPWR VPWR _22940_/A sky130_fd_sc_hd__buf_2
XFILLER_194_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24314_ _25543_/CLK _17652_/X HRESETn VGND VGND VPWR VPWR _17531_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19811__A2_N _19806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21526_ _21525_/Y VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__buf_2
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25294_ _24378_/CLK _13726_/X HRESETn VGND VGND VPWR VPWR _11694_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21102__A _15866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13546__B1 _13481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24245_ _24240_/CLK _24245_/D HRESETn VGND VGND VPWR VPWR _22707_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21608__B2 _21607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21457_ _11728_/X VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__buf_2
XANTENNA__23020__C _23013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12190_ _22285_/A VGND VGND VPWR VPWR _12190_/Y sky130_fd_sc_hd__inv_2
X_20408_ _20408_/A VGND VGND VPWR VPWR _20408_/X sky130_fd_sc_hd__buf_2
X_21388_ _13547_/Y _18277_/X _17455_/X VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__o21a_4
X_24176_ _24192_/CLK _24176_/D HRESETn VGND VGND VPWR VPWR _18474_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23000__A1_N _17322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23127_ _23127_/A VGND VGND VPWR VPWR _23127_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20339_ _21492_/B _20336_/X _20010_/X _20336_/X VGND VGND VPWR VPWR _23429_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21756__B _22575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_76_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_76_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23029__A _22836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23058_ _21314_/A VGND VGND VPWR VPWR _23058_/X sky130_fd_sc_hd__buf_2
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24877__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14900_ _15195_/A VGND VGND VPWR VPWR _15196_/A sky130_fd_sc_hd__inv_2
XANTENNA__22584__A2 _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22009_ _22009_/A _21995_/B VGND VGND VPWR VPWR _22009_/X sky130_fd_sc_hd__and2_4
X_15880_ _15880_/A VGND VGND VPWR VPWR _15880_/X sky130_fd_sc_hd__buf_2
XANTENNA__22868__A _22810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24806__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ _24006_/Q VGND VGND VPWR VPWR _14832_/A sky130_fd_sc_hd__buf_2
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17550_ _11853_/Y _24300_/Q _25553_/Q _17569_/A VGND VGND VPWR VPWR _17555_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14762_ _14759_/X VGND VGND VPWR VPWR _14762_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11974_ _13208_/A VGND VGND VPWR VPWR _11974_/X sky130_fd_sc_hd__buf_2
X_16501_ _16499_/Y _16495_/X _16414_/X _16500_/X VGND VGND VPWR VPWR _24571_/D sky130_fd_sc_hd__a2bb2o_4
X_13713_ _13708_/X _13689_/X _13711_/Y _13712_/X _11705_/A VGND VGND VPWR VPWR _13713_/X
+ sky130_fd_sc_hd__a32o_4
X_17481_ _17480_/X VGND VGND VPWR VPWR _17481_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14693_ _14693_/A VGND VGND VPWR VPWR _14693_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14386__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13290__A _13451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16432_ _16432_/A VGND VGND VPWR VPWR _16432_/Y sky130_fd_sc_hd__inv_2
X_19220_ _19085_/A VGND VGND VPWR VPWR _19220_/X sky130_fd_sc_hd__buf_2
XANTENNA__11803__A _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _13644_/A _14679_/B VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__or2_4
XFILLER_158_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19151_ _19151_/A VGND VGND VPWR VPWR _19151_/X sky130_fd_sc_hd__buf_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _21870_/A VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__inv_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13575_/A VGND VGND VPWR VPWR _13575_/Y sky130_fd_sc_hd__inv_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18102_ _18102_/A VGND VGND VPWR VPWR _18169_/A sky130_fd_sc_hd__buf_2
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15314_ _15142_/Y _15137_/Y _15314_/C VGND VGND VPWR VPWR _15314_/X sky130_fd_sc_hd__or3_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _25431_/Q VGND VGND VPWR VPWR _12616_/A sky130_fd_sc_hd__inv_2
X_19082_ _19090_/A VGND VGND VPWR VPWR _19082_/X sky130_fd_sc_hd__buf_2
X_16294_ HWDATA[30] VGND VGND VPWR VPWR _16294_/X sky130_fd_sc_hd__buf_2
XFILLER_9_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18033_ _13613_/A VGND VGND VPWR VPWR _18037_/A sky130_fd_sc_hd__buf_2
X_15245_ _15053_/X _15218_/X _15208_/X _15241_/Y VGND VGND VPWR VPWR _15245_/X sky130_fd_sc_hd__a211o_4
X_12457_ _12255_/A _12457_/B VGND VGND VPWR VPWR _12457_/X sky130_fd_sc_hd__or2_4
XFILLER_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15176_ _15176_/A VGND VGND VPWR VPWR _15176_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12388_ _12386_/Y _24831_/Q _12387_/X _24828_/Q VGND VGND VPWR VPWR _12388_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14127_ _14126_/X VGND VGND VPWR VPWR _14128_/B sky130_fd_sc_hd__inv_2
X_19984_ _21210_/B _19979_/X _19900_/X _19979_/A VGND VGND VPWR VPWR _23557_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14058_ _14058_/A _14056_/Y _14058_/C _14058_/D VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__and4_4
X_18935_ _18933_/Y _18929_/X _18934_/X _18916_/Y VGND VGND VPWR VPWR _23925_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13009_ _13026_/A _13008_/X VGND VGND VPWR VPWR _13021_/D sky130_fd_sc_hd__or2_4
X_18866_ _18862_/X _18863_/X _18864_/X _18865_/X VGND VGND VPWR VPWR _18872_/C sky130_fd_sc_hd__or4_4
XANTENNA__24547__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17817_ _17896_/A VGND VGND VPWR VPWR _17852_/A sky130_fd_sc_hd__buf_2
XFILLER_94_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ _18797_/A _18795_/A VGND VGND VPWR VPWR _18797_/X sky130_fd_sc_hd__or2_4
XANTENNA__19152__A _19159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17748_ _17896_/A VGND VGND VPWR VPWR _17748_/X sky130_fd_sc_hd__buf_2
XFILLER_36_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17679_ _17585_/D _17678_/X VGND VGND VPWR VPWR _17683_/B sky130_fd_sc_hd__or2_4
XANTENNA__18991__A _19131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19418_ _19148_/A VGND VGND VPWR VPWR _19418_/X sky130_fd_sc_hd__buf_2
X_20690_ _20493_/X _20511_/C _20621_/B VGND VGND VPWR VPWR _24007_/D sky130_fd_sc_hd__o21a_4
XANTENNA__23288__B1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19349_ _19345_/Y _19348_/X _19326_/X _19348_/X VGND VGND VPWR VPWR _23780_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22360_ _21947_/A _22360_/B VGND VGND VPWR VPWR _22362_/B sky130_fd_sc_hd__or2_4
XFILLER_248_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16714__B1 _16534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21311_ _21311_/A VGND VGND VPWR VPWR _21312_/B sky130_fd_sc_hd__buf_2
X_22291_ _24623_/Q _22291_/B VGND VGND VPWR VPWR _22291_/X sky130_fd_sc_hd__or2_4
XFILLER_248_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21242_ _21248_/A VGND VGND VPWR VPWR _21267_/A sky130_fd_sc_hd__buf_2
X_24030_ _24495_/CLK _20766_/X HRESETn VGND VGND VPWR VPWR _13142_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21173_ _15388_/A _21173_/B _21173_/C VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__and3_4
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20124_ _23509_/Q VGND VGND VPWR VPWR _20124_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20055_ _23533_/Q VGND VGND VPWR VPWR _20055_/Y sky130_fd_sc_hd__inv_2
X_24932_ _24354_/CLK _15548_/X HRESETn VGND VGND VPWR VPWR _12073_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_98_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22971__C1 _22970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24863_ _24872_/CLK _15778_/X HRESETn VGND VGND VPWR VPWR _24863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22318__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23814_ _23454_/CLK _23814_/D VGND VGND VPWR VPWR _13413_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24794_ _24794_/CLK _15914_/X HRESETn VGND VGND VPWR VPWR _24794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23669_/CLK _19447_/X VGND VGND VPWR VPWR _18081_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13822__B _13822_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _20956_/Y _20952_/Y VGND VGND VPWR VPWR _20957_/X sky130_fd_sc_hd__and2_4
XPHY_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23279__B1 _12337_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11688_/A _24241_/Q _11688_/Y _22550_/A VGND VGND VPWR VPWR _11697_/B sky130_fd_sc_hd__o22a_4
X_23676_ _24214_/CLK _19654_/X VGND VGND VPWR VPWR _23676_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _13671_/X VGND VGND VPWR VPWR _20888_/Y sky130_fd_sc_hd__inv_2
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25415_ _24867_/CLK _25415_/D HRESETn VGND VGND VPWR VPWR _12557_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22854__C _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22627_ _16776_/A _22543_/X _22544_/X VGND VGND VPWR VPWR _22627_/X sky130_fd_sc_hd__o21a_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ _13456_/A _13352_/X _13360_/C VGND VGND VPWR VPWR _13360_/X sky130_fd_sc_hd__and3_4
X_25346_ _25368_/CLK _13109_/X HRESETn VGND VGND VPWR VPWR _25346_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22558_ _22558_/A VGND VGND VPWR VPWR _23303_/B sky130_fd_sc_hd__buf_2
XFILLER_158_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16705__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12311_ _25356_/Q VGND VGND VPWR VPWR _12311_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13519__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21509_ _21509_/A _21500_/X _21508_/X VGND VGND VPWR VPWR _21509_/X sky130_fd_sc_hd__or3_4
XANTENNA__25005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13291_ _13249_/A _23794_/Q VGND VGND VPWR VPWR _13293_/B sky130_fd_sc_hd__or2_4
X_25277_ _23647_/CLK _25277_/D HRESETn VGND VGND VPWR VPWR _25277_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22489_ _23053_/A VGND VGND VPWR VPWR _22985_/B sky130_fd_sc_hd__buf_2
X_15030_ _15030_/A _15030_/B _15027_/X _15029_/X VGND VGND VPWR VPWR _15031_/D sky130_fd_sc_hd__or4_4
X_12242_ _25439_/Q _12240_/Y _12503_/A _12241_/Y VGND VGND VPWR VPWR _12242_/X sky130_fd_sc_hd__a2bb2o_4
X_24228_ _24230_/CLK _24228_/D HRESETn VGND VGND VPWR VPWR _18273_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14192__B1 _14191_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15765__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _18377_/A _12168_/X _12172_/X VGND VGND VPWR VPWR _12173_/X sky130_fd_sc_hd__a21o_4
X_24159_ _24160_/CLK _18723_/Y HRESETn VGND VGND VPWR VPWR _24159_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16981_ _24397_/Q VGND VGND VPWR VPWR _16981_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18720_ _18720_/A _18720_/B VGND VGND VPWR VPWR _18720_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_100_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24787_/CLK sky130_fd_sc_hd__clkbuf_1
X_15932_ _15655_/X _15844_/X _15851_/X _21023_/B _15931_/X VGND VGND VPWR VPWR _15932_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24640__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_163_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23889_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_6_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15863_ _22684_/B VGND VGND VPWR VPWR _15863_/X sky130_fd_sc_hd__buf_2
X_18651_ _16596_/Y _24145_/Q _16596_/Y _24145_/Q VGND VGND VPWR VPWR _18651_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14814_ _25061_/Q VGND VGND VPWR VPWR _14815_/C sky130_fd_sc_hd__inv_2
X_17602_ _17601_/X VGND VGND VPWR VPWR _24326_/D sky130_fd_sc_hd__inv_2
XFILLER_92_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15794_ _15793_/X VGND VGND VPWR VPWR _15934_/B sky130_fd_sc_hd__buf_2
X_18582_ _18418_/Y _18569_/X VGND VGND VPWR VPWR _18582_/Y sky130_fd_sc_hd__nand2_4
X_14745_ _14744_/X VGND VGND VPWR VPWR _14745_/Y sky130_fd_sc_hd__inv_2
X_17533_ _17526_/X _17533_/B _17533_/C _17532_/X VGND VGND VPWR VPWR _17533_/X sky130_fd_sc_hd__or4_4
X_11957_ _19639_/A VGND VGND VPWR VPWR _11957_/X sky130_fd_sc_hd__buf_2
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17464_ _17464_/A VGND VGND VPWR VPWR _17464_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14676_ _13611_/A _19054_/C _14798_/A VGND VGND VPWR VPWR _14676_/X sky130_fd_sc_hd__o21a_4
X_11888_ _11889_/A _11887_/Y VGND VGND VPWR VPWR _17711_/D sky130_fd_sc_hd__or2_4
X_16415_ _16415_/A VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__buf_2
X_19203_ _19196_/A VGND VGND VPWR VPWR _19203_/X sky130_fd_sc_hd__buf_2
X_13627_ _25076_/Q VGND VGND VPWR VPWR _13628_/B sky130_fd_sc_hd__inv_2
X_17395_ _24000_/Q VGND VGND VPWR VPWR _17396_/A sky130_fd_sc_hd__inv_2
XANTENNA__18316__A _22271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16346_ _16352_/A VGND VGND VPWR VPWR _16346_/X sky130_fd_sc_hd__buf_2
X_19134_ _19134_/A VGND VGND VPWR VPWR _19134_/X sky130_fd_sc_hd__buf_2
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13558_ _25264_/Q VGND VGND VPWR VPWR _13558_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12509_ _12273_/X _12508_/X _12403_/X VGND VGND VPWR VPWR _12509_/Y sky130_fd_sc_hd__a21oi_4
X_19065_ _19065_/A VGND VGND VPWR VPWR _19065_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16277_ _16275_/Y _16196_/X _16276_/X _16196_/X VGND VGND VPWR VPWR _24653_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13489_ _13488_/Y _13486_/X _11847_/X _13486_/X VGND VGND VPWR VPWR _25328_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15228_ _14921_/X _15232_/A _15231_/A _15219_/X VGND VGND VPWR VPWR _15228_/X sky130_fd_sc_hd__or4_4
X_18016_ _18016_/A _18016_/B _18016_/C VGND VGND VPWR VPWR _18028_/B sky130_fd_sc_hd__or3_4
XANTENNA__21677__A _21485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24799__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15675__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15159_ _25001_/Q VGND VGND VPWR VPWR _15362_/A sky130_fd_sc_hd__inv_2
XFILLER_5_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18051__A _18051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24728__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19967_ _19979_/A VGND VGND VPWR VPWR _19967_/X sky130_fd_sc_hd__buf_2
XFILLER_68_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18918_ _18912_/Y _18917_/X _16872_/X _18917_/X VGND VGND VPWR VPWR _18918_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19898_ _21474_/B _19895_/X _19646_/X _19895_/X VGND VGND VPWR VPWR _23590_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18849_ _24565_/Q _18782_/A _16515_/Y _18699_/A VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22301__A _21604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21860_ _14430_/Y _14232_/A _14453_/Y _22334_/B VGND VGND VPWR VPWR _21860_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21508__B1 _18306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20811_ _20808_/Y _20809_/Y _20810_/X VGND VGND VPWR VPWR _20811_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13642__B _13610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21791_ _21648_/A _21791_/B VGND VGND VPWR VPWR _21792_/C sky130_fd_sc_hd__or2_4
XANTENNA__18927__A2_N _18922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23530_ _23514_/CLK _20066_/X VGND VGND VPWR VPWR _20064_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20742_ _20694_/A VGND VGND VPWR VPWR _20765_/A sky130_fd_sc_hd__inv_2
XANTENNA__25516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _23466_/CLK _23461_/D VGND VGND VPWR VPWR _20253_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20673_ _17408_/B VGND VGND VPWR VPWR _20673_/Y sky130_fd_sc_hd__inv_2
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14754__A _14753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25200_ _25200_/CLK _14249_/X HRESETn VGND VGND VPWR VPWR _25200_/Q sky130_fd_sc_hd__dfstp_4
X_22412_ _22854_/B VGND VGND VPWR VPWR _23027_/B sky130_fd_sc_hd__buf_2
X_23392_ _23913_/CLK _20428_/X VGND VGND VPWR VPWR _13278_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25131_ _24337_/CLK _14471_/X HRESETn VGND VGND VPWR VPWR _25131_/Q sky130_fd_sc_hd__dfrtp_4
X_22343_ _17727_/A _22343_/B VGND VGND VPWR VPWR _22343_/X sky130_fd_sc_hd__or2_4
XFILLER_148_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25062_ _25062_/CLK _25062_/D HRESETn VGND VGND VPWR VPWR _25062_/Q sky130_fd_sc_hd__dfrtp_4
X_22274_ _22274_/A _22266_/X _22273_/X VGND VGND VPWR VPWR _22274_/X sky130_fd_sc_hd__and3_4
X_24013_ _25106_/CLK _24013_/D HRESETn VGND VGND VPWR VPWR _24013_/Q sky130_fd_sc_hd__dfrtp_4
X_21225_ _21967_/A _21225_/B _21224_/Y VGND VGND VPWR VPWR _21225_/X sky130_fd_sc_hd__or3_4
XANTENNA__17112__B1 _17065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21156_ _17448_/B _21148_/X _12109_/C _21155_/X VGND VGND VPWR VPWR _21156_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18860__B1 _16517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20107_ _20107_/A VGND VGND VPWR VPWR _20107_/Y sky130_fd_sc_hd__inv_2
X_21087_ _21231_/A VGND VGND VPWR VPWR _22968_/B sky130_fd_sc_hd__buf_2
XFILLER_144_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20038_ _20038_/A VGND VGND VPWR VPWR _20038_/Y sky130_fd_sc_hd__inv_2
X_24915_ _24915_/CLK _24915_/D HRESETn VGND VGND VPWR VPWR _24915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_236_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _23991_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12860_ _12815_/A _12807_/Y _12858_/X _12859_/X VGND VGND VPWR VPWR _12860_/X sky130_fd_sc_hd__or4_4
X_24846_ _24878_/CLK _15819_/X HRESETn VGND VGND VPWR VPWR _12317_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17305__A _17305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23026__B _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20970__B2 _15694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A VGND VGND VPWR VPWR _11811_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11839__A1_N _11837_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _24819_/Q VGND VGND VPWR VPWR _12791_/Y sky130_fd_sc_hd__inv_2
X_24777_ _24777_/CLK _24777_/D HRESETn VGND VGND VPWR VPWR _24777_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _21974_/A _21989_/B VGND VGND VPWR VPWR _21989_/Y sky130_fd_sc_hd__nand2_4
XPHY_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _23969_/Q VGND VGND VPWR VPWR _14530_/X sky130_fd_sc_hd__buf_2
XPHY_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _14417_/A _21045_/A VGND VGND VPWR VPWR _15563_/A sky130_fd_sc_hd__or2_4
X_23728_ _23407_/CLK _23728_/D VGND VGND VPWR VPWR _19493_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16926__B1 _16102_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14116_/A VGND VGND VPWR VPWR _20608_/A sky130_fd_sc_hd__buf_2
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A VGND VGND VPWR VPWR _22745_/A sky130_fd_sc_hd__inv_2
X_23659_ _23642_/CLK _23659_/D VGND VGND VPWR VPWR _23659_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16199_/Y _16197_/X _11755_/X _16197_/X VGND VGND VPWR VPWR _24682_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13412_/A _13412_/B _13411_/X VGND VGND VPWR VPWR _13416_/B sky130_fd_sc_hd__and3_4
X_17180_ _16308_/Y _24371_/Q _16308_/Y _24371_/Q VGND VGND VPWR VPWR _17180_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _14392_/A VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__buf_2
XANTENNA__22475__B2 _22289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16131_ _16130_/Y _16128_/X _15970_/X _16128_/X VGND VGND VPWR VPWR _16131_/X sky130_fd_sc_hd__a2bb2o_4
X_13343_ _13209_/X _13324_/X _13342_/X _25336_/Q _11974_/X VGND VGND VPWR VPWR _13343_/X
+ sky130_fd_sc_hd__o32a_4
X_25329_ _24112_/CLK _13487_/X HRESETn VGND VGND VPWR VPWR _25329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17351__B1 _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16062_ _16060_/Y _16056_/X _15765_/X _16061_/X VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_182_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13274_ _13420_/A _13274_/B VGND VGND VPWR VPWR _13274_/X sky130_fd_sc_hd__or2_4
XFILLER_170_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24892__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15013_ _25029_/Q _15012_/A _15231_/A _15012_/Y VGND VGND VPWR VPWR _15013_/X sky130_fd_sc_hd__o22a_4
XFILLER_185_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20238__B1 _19769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12225_ _25467_/Q VGND VGND VPWR VPWR _12225_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14704__A1_N _21630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12912__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24821__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22105__B _22102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19821_ _19821_/A VGND VGND VPWR VPWR _19821_/Y sky130_fd_sc_hd__inv_2
X_12156_ _24118_/Q _12138_/A VGND VGND VPWR VPWR _12157_/A sky130_fd_sc_hd__and2_4
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17001__A1_N _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_46_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19752_ _13369_/B VGND VGND VPWR VPWR _19752_/Y sky130_fd_sc_hd__inv_2
X_12087_ _12087_/A VGND VGND VPWR VPWR _12087_/Y sky130_fd_sc_hd__inv_2
X_16964_ _16963_/Y VGND VGND VPWR VPWR _16964_/X sky130_fd_sc_hd__buf_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18703_ _18703_/A _18702_/X VGND VGND VPWR VPWR _18711_/A sky130_fd_sc_hd__or2_4
XFILLER_237_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15915_ _15714_/X _15902_/X _15777_/X _21712_/A _15871_/X VGND VGND VPWR VPWR _15915_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_204_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19683_ _19681_/Y _19676_/X _19659_/X _19682_/X VGND VGND VPWR VPWR _23666_/D sky130_fd_sc_hd__a2bb2o_4
X_16895_ _16893_/Y _16889_/X _16894_/X _16889_/X VGND VGND VPWR VPWR _16895_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22121__A _22121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18634_ _24539_/Q _24150_/Q _16583_/Y _18698_/C VGND VGND VPWR VPWR _18642_/A sky130_fd_sc_hd__o22a_4
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15846_ _15833_/X _15844_/X _15777_/X _24828_/Q _15802_/A VGND VGND VPWR VPWR _15846_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15661__C _15661_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18565_ _18515_/A _18565_/B VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__or2_4
X_12989_ _12989_/A VGND VGND VPWR VPWR _12989_/Y sky130_fd_sc_hd__inv_2
X_15777_ _11861_/A VGND VGND VPWR VPWR _15777_/X sky130_fd_sc_hd__buf_2
XFILLER_18_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22163__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16272__A1_N _16271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_HCLK clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _24315_/Q VGND VGND VPWR VPWR _17516_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14728_ _14728_/A _14728_/B _14722_/X _14727_/X VGND VGND VPWR VPWR _14729_/A sky130_fd_sc_hd__or4_4
X_18496_ _18496_/A VGND VGND VPWR VPWR _18496_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16917__B1 _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14659_ _17985_/A VGND VGND VPWR VPWR _18013_/A sky130_fd_sc_hd__buf_2
X_17447_ _21020_/A VGND VGND VPWR VPWR _17447_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18046__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22466__A1 _16259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17378_ _17378_/A _17378_/B VGND VGND VPWR VPWR _17378_/Y sky130_fd_sc_hd__nand2_4
XFILLER_220_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19117_ _19116_/Y _19112_/X _18934_/X _19099_/Y VGND VGND VPWR VPWR _19117_/X sky130_fd_sc_hd__a2bb2o_4
X_16329_ _24634_/Q VGND VGND VPWR VPWR _16329_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24909__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19048_ _19048_/A VGND VGND VPWR VPWR _19048_/X sky130_fd_sc_hd__buf_2
XFILLER_161_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24562__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21010_ _21010_/A _24343_/Q VGND VGND VPWR VPWR _21010_/X sky130_fd_sc_hd__and2_4
XFILLER_114_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21854__B _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22961_ _12834_/Y _21456_/X _16950_/Y _22839_/X VGND VGND VPWR VPWR _22961_/X sky130_fd_sc_hd__o22a_4
X_24700_ _24689_/CLK _24700_/D HRESETn VGND VGND VPWR VPWR _16140_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20401__B1 _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21912_ _21907_/X _21911_/X _22221_/A VGND VGND VPWR VPWR _21912_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18070__A1 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22892_ _22801_/X _22890_/X _22804_/X _22891_/X VGND VGND VPWR VPWR _22893_/B sky130_fd_sc_hd__o22a_4
XFILLER_244_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21292__D _21291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16081__B1 _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24631_ _24629_/CLK _16340_/X HRESETn VGND VGND VPWR VPWR _16338_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21843_ _21842_/Y _21324_/X _24488_/Q _22891_/B VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_66_0_HCLK clkbuf_8_66_0_HCLK/A VGND VGND VPWR VPWR _25444_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_82_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24562_ _24562_/CLK _24562_/D HRESETn VGND VGND VPWR VPWR _16522_/A sky130_fd_sc_hd__dfrtp_4
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21774_ _21629_/A _20138_/Y VGND VGND VPWR VPWR _21775_/C sky130_fd_sc_hd__or2_4
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _23513_/CLK _23513_/D VGND VGND VPWR VPWR _23513_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725_ _20725_/A _20725_/B VGND VGND VPWR VPWR _20725_/X sky130_fd_sc_hd__or2_4
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24493_ _24493_/CLK _16707_/X HRESETn VGND VGND VPWR VPWR _16706_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _24343_/CLK _23444_/D VGND VGND VPWR VPWR _23444_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20656_ _23994_/Q _20653_/A VGND VGND VPWR VPWR _20656_/Y sky130_fd_sc_hd__nand2_4
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17795__A _16910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23375_ _23362_/X VGND VGND VPWR VPWR IRQ[19] sky130_fd_sc_hd__buf_2
X_20587_ _20587_/A VGND VGND VPWR VPWR _23956_/D sky130_fd_sc_hd__inv_2
XFILLER_164_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25114_ _23970_/CLK _14527_/X HRESETn VGND VGND VPWR VPWR _20609_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_192_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22326_ _22326_/A VGND VGND VPWR VPWR _22327_/D sky130_fd_sc_hd__inv_2
XFILLER_125_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25045_ _25023_/CLK _25045_/D HRESETn VGND VGND VPWR VPWR pwm_S6 sky130_fd_sc_hd__dfrtp_4
XFILLER_124_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22257_ _21685_/X _22257_/B _22256_/X VGND VGND VPWR VPWR _22257_/X sky130_fd_sc_hd__and3_4
X_12010_ _12010_/A VGND VGND VPWR VPWR _12010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14650__C _14650_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12173__A2 _12168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21208_ _21211_/A _20033_/Y VGND VGND VPWR VPWR _21208_/X sky130_fd_sc_hd__or2_4
XANTENNA__18833__B1 _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22188_ _21578_/X _22186_/X _21584_/X _22187_/X VGND VGND VPWR VPWR _22188_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21139_ _23939_/Q VGND VGND VPWR VPWR _21139_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13961_ _13958_/A _13950_/Y _13952_/C _13960_/Y VGND VGND VPWR VPWR _14259_/A sky130_fd_sc_hd__and4_4
X_12912_ _12912_/A _12912_/B _12911_/X VGND VGND VPWR VPWR _12921_/D sky130_fd_sc_hd__or3_4
X_15700_ _15699_/X VGND VGND VPWR VPWR _15700_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16680_ _16685_/A VGND VGND VPWR VPWR _16680_/X sky130_fd_sc_hd__buf_2
X_13892_ _24007_/Q _13891_/X _14284_/A _13876_/A VGND VGND VPWR VPWR _13892_/X sky130_fd_sc_hd__o22a_4
XFILLER_219_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21780__A _22090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12843_ _12969_/A _22302_/A _12837_/Y _21712_/A VGND VGND VPWR VPWR _12843_/X sky130_fd_sc_hd__a2bb2o_4
X_15631_ _15631_/A VGND VGND VPWR VPWR _15631_/Y sky130_fd_sc_hd__inv_2
X_24829_ _24825_/CLK _24829_/D HRESETn VGND VGND VPWR VPWR _24829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15562_ HWDATA[31] VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__buf_2
X_18350_ _13183_/X _18352_/A _18347_/X VGND VGND VPWR VPWR _18350_/X sky130_fd_sc_hd__o21a_4
X_12774_ _22875_/A VGND VGND VPWR VPWR _12774_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _25117_/Q _14517_/A _14524_/A _14512_/Y VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__a211o_4
X_17301_ _17266_/A _17300_/X VGND VGND VPWR VPWR _17301_/X sky130_fd_sc_hd__or2_4
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _15791_/C VGND VGND VPWR VPWR _16378_/C sky130_fd_sc_hd__buf_2
XFILLER_203_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15493_/A _15493_/B VGND VGND VPWR VPWR _20437_/A sky130_fd_sc_hd__nor2_4
X_18281_ _24224_/Q VGND VGND VPWR VPWR _19527_/C sky130_fd_sc_hd__buf_2
XFILLER_159_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _22334_/B VGND VGND VPWR VPWR _15471_/A sky130_fd_sc_hd__buf_2
X_17232_ _16317_/A _17231_/Y _16322_/Y _17229_/A VGND VGND VPWR VPWR _17232_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11656_/A VGND VGND VPWR VPWR _11970_/C sky130_fd_sc_hd__buf_2
XANTENNA__21004__B _14205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22448__B2 _21547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17163_ _17053_/C _17136_/X VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__or2_4
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _25162_/Q _14360_/A _25161_/Q _14354_/B VGND VGND VPWR VPWR _14375_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17324__B1 _17288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ _16113_/Y _16111_/X _11773_/X _16111_/X VGND VGND VPWR VPWR _16114_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13326_ _13245_/X _13326_/B VGND VGND VPWR VPWR _13326_/X sky130_fd_sc_hd__or2_4
X_17094_ _24401_/Q _17094_/B VGND VGND VPWR VPWR _17094_/X sky130_fd_sc_hd__or2_4
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15886__B1 _11783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16045_ _16042_/Y _16044_/X _11805_/X _16044_/X VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__a2bb2o_4
X_13257_ _13443_/A VGND VGND VPWR VPWR _13257_/X sky130_fd_sc_hd__buf_2
XFILLER_142_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12208_ _12208_/A VGND VGND VPWR VPWR _12208_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13188_ _13178_/A _23876_/Q VGND VGND VPWR VPWR _13188_/X sky130_fd_sc_hd__or2_4
XFILLER_124_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19804_ _21766_/B _19797_/X _19803_/X _19797_/X VGND VGND VPWR VPWR _23624_/D sky130_fd_sc_hd__a2bb2o_4
X_12139_ _24117_/Q _12150_/A _12138_/Y VGND VGND VPWR VPWR _20982_/A sky130_fd_sc_hd__o21a_4
XANTENNA__15953__A _15947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17996_ _17991_/X _17996_/B _17995_/X VGND VGND VPWR VPWR _17996_/X sky130_fd_sc_hd__and3_4
XFILLER_215_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22908__C1 _22907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19735_ _19732_/Y _19733_/X _19734_/X _19733_/X VGND VGND VPWR VPWR _23647_/D sky130_fd_sc_hd__a2bb2o_4
X_16947_ _16120_/Y _24285_/Q _22574_/A _17861_/C VGND VGND VPWR VPWR _16947_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12368__A2_N _24840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19666_ _13397_/B VGND VGND VPWR VPWR _19666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16878_ _16875_/Y _16868_/X _16876_/X _16877_/X VGND VGND VPWR VPWR _16878_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18617_ _24152_/Q VGND VGND VPWR VPWR _18617_/Y sky130_fd_sc_hd__inv_2
X_15829_ _15825_/X _15828_/X _16238_/A _24840_/Q _15826_/X VGND VGND VPWR VPWR _24840_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_231_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19597_ _21382_/C VGND VGND VPWR VPWR _19597_/X sky130_fd_sc_hd__buf_2
XANTENNA__22136__B1 _22123_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15810__B1 _11763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18548_ _18550_/A _18548_/B _18548_/C VGND VGND VPWR VPWR _24180_/D sky130_fd_sc_hd__and3_4
XFILLER_240_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18479_ _18595_/A _18425_/Y _18479_/C _18479_/D VGND VGND VPWR VPWR _18479_/X sky130_fd_sc_hd__or4_4
XANTENNA__12817__A _12817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20510_ _14286_/Y _20503_/B _24093_/Q VGND VGND VPWR VPWR _20510_/X sky130_fd_sc_hd__and3_4
X_21490_ _21687_/A _21490_/B VGND VGND VPWR VPWR _21490_/X sky130_fd_sc_hd__or2_4
XFILLER_147_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20441_ _14395_/A _23938_/D _20463_/C VGND VGND VPWR VPWR _20442_/A sky130_fd_sc_hd__o21a_4
XANTENNA__24743__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23160_ _23113_/X _23158_/X _23159_/X _24851_/Q _23115_/X VGND VGND VPWR VPWR _23160_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_180_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20372_ _20372_/A VGND VGND VPWR VPWR _20372_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21662__A2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22111_ _23253_/A _22111_/B _22110_/X VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__and3_4
X_23091_ _23091_/A _22954_/B _22830_/C VGND VGND VPWR VPWR _23091_/X sky130_fd_sc_hd__and3_4
X_22042_ _22028_/A _19631_/Y VGND VGND VPWR VPWR _22043_/C sky130_fd_sc_hd__or2_4
XFILLER_142_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15863__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23993_ _23998_/CLK _20655_/Y HRESETn VGND VGND VPWR VPWR _17402_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14479__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22944_ _22944_/A _22939_/X _22944_/C VGND VGND VPWR VPWR _22944_/X sky130_fd_sc_hd__and3_4
XANTENNA__25531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16054__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22875_ _22875_/A _22985_/B VGND VGND VPWR VPWR _22875_/X sky130_fd_sc_hd__or2_4
XFILLER_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14629__D _13547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24614_ _25011_/CLK _16392_/X HRESETn VGND VGND VPWR VPWR _24614_/Q sky130_fd_sc_hd__dfrtp_4
X_21826_ _21497_/A _21826_/B VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__or2_4
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24545_ _24562_/CLK _24545_/D HRESETn VGND VGND VPWR VPWR _24545_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21757_ _21757_/A _21330_/A VGND VGND VPWR VPWR _21757_/X sky130_fd_sc_hd__and2_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17554__B1 _11789_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23023__C _22954_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _24018_/Q VGND VGND VPWR VPWR _20708_/Y sky130_fd_sc_hd__inv_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12489_/X VGND VGND VPWR VPWR _12491_/B sky130_fd_sc_hd__inv_2
X_24476_ _24476_/CLK _16751_/X HRESETn VGND VGND VPWR VPWR _16750_/A sky130_fd_sc_hd__dfrtp_4
X_21688_ _21688_/A _21688_/B VGND VGND VPWR VPWR _21689_/C sky130_fd_sc_hd__or2_4
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23427_ _23493_/CLK _23427_/D VGND VGND VPWR VPWR _21996_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20639_ _17399_/X _20639_/B _20628_/X VGND VGND VPWR VPWR _20639_/X sky130_fd_sc_hd__and3_4
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _14138_/X _14159_/X _25143_/Q _14145_/X VGND VGND VPWR VPWR _14160_/Y sky130_fd_sc_hd__a22oi_4
X_23358_ _23358_/A _23358_/B VGND VGND VPWR VPWR _23358_/Y sky130_fd_sc_hd__nor2_4
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16747__A1_N _15024_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13111_ _12351_/A _13111_/B VGND VGND VPWR VPWR _13111_/X sky130_fd_sc_hd__or2_4
X_22309_ _12842_/A _22306_/X _22308_/X VGND VGND VPWR VPWR _22309_/X sky130_fd_sc_hd__a21o_4
XANTENNA__19059__B1 _19008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14091_ _14027_/A _14090_/X _14087_/X _13999_/D _14085_/X VGND VGND VPWR VPWR _14091_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23289_ _23321_/A _23288_/X VGND VGND VPWR VPWR _23289_/X sky130_fd_sc_hd__and2_4
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_222_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13042_ _12308_/Y _13044_/B _13041_/Y VGND VGND VPWR VPWR _13042_/X sky130_fd_sc_hd__o21a_4
X_25028_ _25023_/CLK _25028_/D HRESETn VGND VGND VPWR VPWR _14969_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21775__A _21630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15883__A3 _15734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17850_ _17762_/A _17849_/Y VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__or2_4
X_16801_ _24451_/Q VGND VGND VPWR VPWR _16801_/Y sky130_fd_sc_hd__inv_2
X_17781_ _17773_/X _17780_/X VGND VGND VPWR VPWR _17781_/X sky130_fd_sc_hd__or2_4
X_14993_ _14993_/A _14993_/B _14983_/X _14992_/X VGND VGND VPWR VPWR _14994_/B sky130_fd_sc_hd__or4_4
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19520_ _19507_/Y VGND VGND VPWR VPWR _19520_/X sky130_fd_sc_hd__buf_2
XANTENNA__22905__A2 _22541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16732_ _16731_/Y VGND VGND VPWR VPWR _16733_/A sky130_fd_sc_hd__buf_2
XANTENNA__19231__B1 _19139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13944_ _13944_/A _13941_/Y _13933_/X _13943_/X VGND VGND VPWR VPWR _13945_/A sky130_fd_sc_hd__or4_4
XANTENNA__25272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20287__A2_N _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16045__B1 _11805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19451_ _19438_/A VGND VGND VPWR VPWR _19451_/X sky130_fd_sc_hd__buf_2
XFILLER_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13875_ _20681_/A _13870_/X _25255_/Q _13872_/X VGND VGND VPWR VPWR _13875_/X sky130_fd_sc_hd__o22a_4
X_16663_ _16662_/Y _16660_/X _16395_/X _16660_/X VGND VGND VPWR VPWR _24511_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18402_ _16212_/Y _24188_/Q _16212_/Y _24188_/Q VGND VGND VPWR VPWR _18402_/X sky130_fd_sc_hd__a2bb2o_4
X_12826_ _12825_/Y _24812_/Q _25383_/Q _12764_/Y VGND VGND VPWR VPWR _12836_/A sky130_fd_sc_hd__a2bb2o_4
X_15614_ _15614_/A VGND VGND VPWR VPWR _15614_/X sky130_fd_sc_hd__buf_2
XFILLER_234_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19382_ _19368_/Y VGND VGND VPWR VPWR _19382_/X sky130_fd_sc_hd__buf_2
X_16594_ _16594_/A VGND VGND VPWR VPWR _16594_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20210__A2_N _20205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18333_ _18959_/A _18333_/B _18333_/C _19075_/B VGND VGND VPWR VPWR _18333_/X sky130_fd_sc_hd__and4_4
X_12757_ _12842_/A _12755_/Y _12864_/A _23199_/A VGND VGND VPWR VPWR _12760_/C sky130_fd_sc_hd__a2bb2o_4
X_15545_ _12068_/X _15544_/X HADDR[4] _15544_/X VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12637__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11699_/X _11708_/B _11704_/X _11708_/D VGND VGND VPWR VPWR _11708_/X sky130_fd_sc_hd__or4_4
X_15476_ _24961_/Q VGND VGND VPWR VPWR _15476_/Y sky130_fd_sc_hd__inv_2
X_18264_ _11703_/Y _18258_/X _16861_/X _18243_/A VGND VGND VPWR VPWR _24233_/D sky130_fd_sc_hd__a2bb2o_4
X_12688_ _12618_/B _12685_/D VGND VGND VPWR VPWR _12689_/B sky130_fd_sc_hd__or2_4
XFILLER_147_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20854__A _20854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15020__B2 _15019_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _14427_/A VGND VGND VPWR VPWR _14427_/X sky130_fd_sc_hd__buf_2
X_17215_ _17214_/Y VGND VGND VPWR VPWR _17391_/A sky130_fd_sc_hd__buf_2
XFILLER_147_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15948__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18195_ _18131_/A _18191_/X _18195_/C VGND VGND VPWR VPWR _18203_/B sky130_fd_sc_hd__or3_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _14347_/A _14360_/A VGND VGND VPWR VPWR _14358_/X sky130_fd_sc_hd__or2_4
X_17146_ _17050_/C _17144_/X _17145_/Y VGND VGND VPWR VPWR _17146_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _13412_/A _13307_/X _13309_/C VGND VGND VPWR VPWR _13315_/B sky130_fd_sc_hd__and3_4
X_17077_ _17034_/A _17075_/X _17076_/X _17070_/Y VGND VGND VPWR VPWR _17078_/A sky130_fd_sc_hd__a211o_4
X_14289_ _15446_/A VGND VGND VPWR VPWR _14289_/X sky130_fd_sc_hd__buf_2
X_16028_ _16028_/A VGND VGND VPWR VPWR _16028_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15874__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15683__A _16382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17979_ _17979_/A _19394_/A VGND VGND VPWR VPWR _17979_/X sky130_fd_sc_hd__or2_4
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19718_ _17463_/X _20079_/B _20079_/C _18905_/D VGND VGND VPWR VPWR _19719_/A sky130_fd_sc_hd__or4_4
XFILLER_226_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20990_ _24126_/Q _24124_/Q VGND VGND VPWR VPWR _20990_/X sky130_fd_sc_hd__and2_4
XFILLER_226_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19649_ _21195_/B _19642_/X _19501_/X _19624_/Y VGND VGND VPWR VPWR _19649_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15909__A1_N _12778_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22660_ _22660_/A VGND VGND VPWR VPWR _22660_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21611_ _21260_/A VGND VGND VPWR VPWR _21611_/X sky130_fd_sc_hd__buf_2
XFILLER_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22591_ _16845_/A _22541_/X _22542_/X _22590_/X VGND VGND VPWR VPWR _22591_/X sky130_fd_sc_hd__a211o_4
XFILLER_240_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12245__A2_N _22644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24330_ _24194_/CLK _17453_/X HRESETn VGND VGND VPWR VPWR _21020_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21542_ _21542_/A VGND VGND VPWR VPWR _21542_/X sky130_fd_sc_hd__buf_2
XANTENNA__21883__A2 _21881_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24261_ _23597_/CLK _17916_/X HRESETn VGND VGND VPWR VPWR _17900_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_5_16_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15858__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21473_ _21473_/A VGND VGND VPWR VPWR _21474_/A sky130_fd_sc_hd__buf_2
XANTENNA__18234__A _18234_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23212_ _16662_/Y _23303_/B VGND VGND VPWR VPWR _23212_/X sky130_fd_sc_hd__and2_4
X_20424_ _20422_/Y _18907_/X _19817_/X _20423_/X VGND VGND VPWR VPWR _23394_/D sky130_fd_sc_hd__a2bb2o_4
X_24192_ _24192_/CLK _24192_/D HRESETn VGND VGND VPWR VPWR _24192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23143_ _22813_/A VGND VGND VPWR VPWR _23156_/A sky130_fd_sc_hd__buf_2
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20355_ _20342_/X _19599_/D _15993_/X _21995_/B _20346_/X VGND VGND VPWR VPWR _20355_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23074_ _23008_/A _23073_/X VGND VGND VPWR VPWR _23074_/Y sky130_fd_sc_hd__nor2_4
X_20286_ _23449_/Q VGND VGND VPWR VPWR _21921_/B sky130_fd_sc_hd__inv_2
XFILLER_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22596__B1 _21968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22025_ _22036_/A _22025_/B _22025_/C VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__and3_4
XFILLER_0_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24121__D MSI_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22899__A1 _24538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11990_ _11663_/A _11663_/B _11985_/X VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__and3_4
X_23976_ _23976_/CLK _23976_/D HRESETn VGND VGND VPWR VPWR _21369_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16027__B1 _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22927_ _22306_/A VGND VGND VPWR VPWR _22927_/X sky130_fd_sc_hd__buf_2
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13660_ _13660_/A VGND VGND VPWR VPWR _13660_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22858_ _21881_/X VGND VGND VPWR VPWR _22858_/X sky130_fd_sc_hd__buf_2
XFILLER_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_36_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12611_ _12638_/B VGND VGND VPWR VPWR _12730_/A sky130_fd_sc_hd__buf_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21809_ _21805_/X _21808_/X _17732_/X VGND VGND VPWR VPWR _21809_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13591_ _25092_/Q VGND VGND VPWR VPWR _14613_/A sky130_fd_sc_hd__inv_2
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22789_ _24633_/Q _22789_/B VGND VGND VPWR VPWR _22789_/X sky130_fd_sc_hd__or2_4
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_99_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21323__B2 _21322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24665__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15330_ _15329_/X VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__inv_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12542_ _24879_/Q VGND VGND VPWR VPWR _12542_/Y sky130_fd_sc_hd__inv_2
X_24528_ _24528_/CLK _16614_/X HRESETn VGND VGND VPWR VPWR _16612_/A sky130_fd_sc_hd__dfrtp_4
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15261_ _15260_/X VGND VGND VPWR VPWR _15261_/Y sky130_fd_sc_hd__inv_2
X_12473_ _12458_/A _12473_/B _12472_/X VGND VGND VPWR VPWR _25451_/D sky130_fd_sc_hd__and3_4
X_24459_ _25018_/CLK _16784_/X HRESETn VGND VGND VPWR VPWR _15017_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16686__A1_N _16684_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14212_ _20524_/A VGND VGND VPWR VPWR _20518_/A sky130_fd_sc_hd__inv_2
X_17000_ _24395_/Q VGND VGND VPWR VPWR _17118_/A sky130_fd_sc_hd__inv_2
XFILLER_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15192_ _15191_/X VGND VGND VPWR VPWR _15192_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_HCLK clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14143_ _23967_/D _14142_/X _14425_/A _23967_/D VGND VGND VPWR VPWR _14143_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17983__A _18006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14074_ _14082_/A VGND VGND VPWR VPWR _14074_/X sky130_fd_sc_hd__buf_2
X_18951_ _23919_/Q VGND VGND VPWR VPWR _18951_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13025_ _13044_/A _13025_/B _13025_/C VGND VGND VPWR VPWR _13025_/X sky130_fd_sc_hd__and3_4
X_17902_ _17900_/Y _17913_/B _17900_/A _17901_/Y VGND VGND VPWR VPWR _17907_/A sky130_fd_sc_hd__o22a_4
X_18882_ _20579_/A _18881_/X VGND VGND VPWR VPWR _18883_/B sky130_fd_sc_hd__or2_4
XANTENNA__25453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17833_ _16914_/Y _17832_/X VGND VGND VPWR VPWR _17833_/Y sky130_fd_sc_hd__nand2_4
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22339__B1 _14227_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15653__D _14442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19204__B1 _19091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ _17764_/A VGND VGND VPWR VPWR _17766_/A sky130_fd_sc_hd__inv_2
XANTENNA__16281__A3 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14976_ _14976_/A VGND VGND VPWR VPWR _14976_/Y sky130_fd_sc_hd__inv_2
X_19503_ _23724_/Q VGND VGND VPWR VPWR _22343_/B sky130_fd_sc_hd__inv_2
XFILLER_207_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16715_ _24489_/Q VGND VGND VPWR VPWR _16715_/Y sky130_fd_sc_hd__inv_2
X_13927_ _13927_/A _13927_/B _13927_/C _13903_/Y VGND VGND VPWR VPWR _13927_/X sky130_fd_sc_hd__and4_4
X_17695_ _17674_/X _17695_/B _17702_/C VGND VGND VPWR VPWR _24301_/D sky130_fd_sc_hd__and3_4
XFILLER_207_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19434_ _19433_/Y _19429_/X _19410_/X _19415_/A VGND VGND VPWR VPWR _23749_/D sky130_fd_sc_hd__a2bb2o_4
X_16646_ _16646_/A VGND VGND VPWR VPWR _24517_/D sky130_fd_sc_hd__inv_2
X_13858_ _13857_/Y _13838_/A _13819_/X _13838_/A VGND VGND VPWR VPWR _25260_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _12941_/A _22641_/A _12807_/Y _22641_/A VGND VGND VPWR VPWR _12809_/X sky130_fd_sc_hd__a2bb2o_4
X_19365_ _19364_/Y _19360_/X _19254_/X _19353_/A VGND VGND VPWR VPWR _19365_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16577_ _16576_/Y _16572_/X _16407_/X _16572_/X VGND VGND VPWR VPWR _24542_/D sky130_fd_sc_hd__a2bb2o_4
X_13789_ _13789_/A VGND VGND VPWR VPWR _13789_/X sky130_fd_sc_hd__buf_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18715__C1 _18714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18316_ _22271_/A VGND VGND VPWR VPWR _21676_/A sky130_fd_sc_hd__buf_2
XANTENNA__22454__A1_N _17861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14979__A2_N _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15528_ _11739_/A VGND VGND VPWR VPWR _15528_/Y sky130_fd_sc_hd__inv_2
X_19296_ _19295_/Y _19293_/X _16897_/X _19293_/X VGND VGND VPWR VPWR _23798_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21865__A2 _12107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20164__A2_N _20163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18247_ _20408_/A VGND VGND VPWR VPWR _18247_/X sky130_fd_sc_hd__buf_2
XANTENNA__15678__A _21596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15459_ _13963_/A _15458_/X _15455_/X _13952_/C _15453_/X VGND VGND VPWR VPWR _24972_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18178_ _18178_/A _18178_/B VGND VGND VPWR VPWR _18178_/X sky130_fd_sc_hd__or2_4
XFILLER_144_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17129_ _17129_/A _17129_/B VGND VGND VPWR VPWR _17132_/B sky130_fd_sc_hd__or2_4
XANTENNA__17893__A _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20140_ _20140_/A VGND VGND VPWR VPWR _21629_/B sky130_fd_sc_hd__inv_2
XFILLER_143_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20071_ _20071_/A VGND VGND VPWR VPWR _20071_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23830_ _23830_/CLK _23830_/D VGND VGND VPWR VPWR _19205_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22958__B _23027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16009__B1 _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23761_ _23768_/CLK _19400_/X VGND VGND VPWR VPWR _18074_/B sky130_fd_sc_hd__dfxtp_4
X_20973_ _12015_/A _20972_/B VGND VGND VPWR VPWR _20973_/X sky130_fd_sc_hd__and2_4
X_22712_ _16427_/A _22316_/B VGND VGND VPWR VPWR _22715_/B sky130_fd_sc_hd__or2_4
X_25500_ _24201_/CLK _12039_/X HRESETn VGND VGND VPWR VPWR _25500_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23692_ _23400_/CLK _19602_/X VGND VGND VPWR VPWR _23692_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25431_ _25425_/CLK _25431_/D HRESETn VGND VGND VPWR VPWR _25431_/Q sky130_fd_sc_hd__dfrtp_4
X_22643_ _21060_/A _22643_/B VGND VGND VPWR VPWR _22643_/Y sky130_fd_sc_hd__nand2_4
XFILLER_198_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15783__A2 _15774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25362_ _25358_/CLK _25362_/D HRESETn VGND VGND VPWR VPWR _12370_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22574_ _22574_/A _21103_/A VGND VGND VPWR VPWR _22574_/X sky130_fd_sc_hd__or2_4
XANTENNA__21856__A2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24313_ _25543_/CLK _24313_/D HRESETn VGND VGND VPWR VPWR _17535_/A sky130_fd_sc_hd__dfrtp_4
X_21525_ _21967_/A VGND VGND VPWR VPWR _21525_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25293_ _25292_/CLK _13728_/X HRESETn VGND VGND VPWR VPWR _11676_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_194_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24244_ _24240_/CLK _24244_/D HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21456_ _21027_/X VGND VGND VPWR VPWR _21456_/X sky130_fd_sc_hd__buf_2
XFILLER_181_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20407_ _20342_/X _20404_/X _13844_/A _22408_/A _20406_/X VGND VGND VPWR VPWR _23403_/D
+ sky130_fd_sc_hd__a32o_4
X_24175_ _24192_/CLK _24175_/D HRESETn VGND VGND VPWR VPWR _18475_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21387_ _21974_/A _21385_/X _13792_/A _21386_/X VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__a211o_4
XFILLER_134_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16496__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23126_ _23124_/X _23125_/X _23058_/X _16021_/A _22990_/X VGND VGND VPWR VPWR _23127_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20292__B2 _20291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20338_ _20338_/A VGND VGND VPWR VPWR _21492_/B sky130_fd_sc_hd__inv_2
XANTENNA__12752__A2_N _22605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18237__A1 _17973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23057_ _16314_/A _23165_/B VGND VGND VPWR VPWR _23057_/X sky130_fd_sc_hd__or2_4
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19434__B1 _19410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20269_ _23455_/Q VGND VGND VPWR VPWR _20269_/Y sky130_fd_sc_hd__inv_2
X_22008_ _17900_/Y _23422_/Q _22009_/A _21995_/B VGND VGND VPWR VPWR _22008_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14830_ _14227_/A _14819_/X _14820_/X _14829_/Y VGND VGND VPWR VPWR _14830_/X sky130_fd_sc_hd__o22a_4
XFILLER_248_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11973_ _11973_/A VGND VGND VPWR VPWR _13208_/A sky130_fd_sc_hd__buf_2
X_14761_ _14761_/A _14753_/X VGND VGND VPWR VPWR _14761_/X sky130_fd_sc_hd__and2_4
XFILLER_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23959_ _23960_/CLK _20599_/Y HRESETn VGND VGND VPWR VPWR _23959_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13482__B1 _13481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24846__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _16495_/A VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__buf_2
XFILLER_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13712_ _13686_/Y VGND VGND VPWR VPWR _13712_/X sky130_fd_sc_hd__buf_2
X_14692_ _14692_/A _14692_/B VGND VGND VPWR VPWR _14693_/A sky130_fd_sc_hd__and2_4
X_17480_ _13200_/A _17479_/Y _13200_/A _17479_/Y VGND VGND VPWR VPWR _17480_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14386__B _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16420__B1 _16419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16431_ _16430_/Y _16428_/X _16245_/X _16428_/X VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13643_ _13643_/A VGND VGND VPWR VPWR _13644_/A sky130_fd_sc_hd__inv_2
XFILLER_232_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23297__A1 _22563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25075__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19150_ _19150_/A VGND VGND VPWR VPWR _19150_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13574_ _25262_/Q VGND VGND VPWR VPWR _13574_/Y sky130_fd_sc_hd__inv_2
X_16362_ _16361_/Y _16359_/X _16073_/X _16359_/X VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18101_ _18166_/A _18101_/B _18100_/X VGND VGND VPWR VPWR _18106_/B sky130_fd_sc_hd__and3_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12525_ _25412_/Q _12523_/Y _12642_/B _12536_/A VGND VGND VPWR VPWR _12525_/X sky130_fd_sc_hd__a2bb2o_4
X_15313_ _15308_/X _15310_/X _15312_/X VGND VGND VPWR VPWR _15314_/C sky130_fd_sc_hd__or3_4
XFILLER_9_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15498__A _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16293_ _24647_/Q VGND VGND VPWR VPWR _16293_/Y sky130_fd_sc_hd__inv_2
X_19081_ _13270_/B VGND VGND VPWR VPWR _19081_/Y sky130_fd_sc_hd__inv_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_123_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24503_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_185_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18032_ _17973_/X _18030_/X _24253_/Q _18031_/X VGND VGND VPWR VPWR _18032_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_186_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _23918_/CLK sky130_fd_sc_hd__clkbuf_1
X_12456_ _12453_/B VGND VGND VPWR VPWR _12457_/B sky130_fd_sc_hd__inv_2
X_15244_ _15252_/A _15244_/B _15243_/X VGND VGND VPWR VPWR _25028_/D sky130_fd_sc_hd__and3_4
XFILLER_200_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15175_ _15182_/A _15182_/B _14986_/Y _15174_/X VGND VGND VPWR VPWR _15176_/A sky130_fd_sc_hd__or4_4
X_12387_ _12381_/Y VGND VGND VPWR VPWR _12387_/X sky130_fd_sc_hd__buf_2
XFILLER_125_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14126_ _25226_/Q _14125_/X _14112_/A VGND VGND VPWR VPWR _14126_/X sky130_fd_sc_hd__or3_4
XFILLER_114_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15829__A3 _16238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19983_ _19983_/A VGND VGND VPWR VPWR _21210_/B sky130_fd_sc_hd__inv_2
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14057_ _14057_/A VGND VGND VPWR VPWR _14058_/D sky130_fd_sc_hd__inv_2
X_18934_ _20146_/A VGND VGND VPWR VPWR _18934_/X sky130_fd_sc_hd__buf_2
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19425__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16239__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13008_ _13038_/A _12370_/Y _12995_/X _13007_/X VGND VGND VPWR VPWR _13008_/X sky130_fd_sc_hd__or4_4
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18865_ _24573_/Q _18756_/A _24579_/Q _18703_/A VGND VGND VPWR VPWR _18865_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17816_ _17816_/A VGND VGND VPWR VPWR _17816_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18796_ _18604_/X _18795_/Y VGND VGND VPWR VPWR _18796_/X sky130_fd_sc_hd__or2_4
XFILLER_36_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17747_ _16962_/X VGND VGND VPWR VPWR _17896_/A sky130_fd_sc_hd__buf_2
X_14959_ _14958_/Y _24433_/Q _14958_/Y _24433_/Q VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18049__A _18234_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24587__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13481__A _13481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17678_ _17684_/A _17684_/B VGND VGND VPWR VPWR _17678_/X sky130_fd_sc_hd__or2_4
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16411__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19417_ _23755_/Q VGND VGND VPWR VPWR _19417_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16629_ _24521_/Q VGND VGND VPWR VPWR _16629_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16792__A _16737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12830__A1_N _12828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19348_ _19353_/A VGND VGND VPWR VPWR _19348_/X sky130_fd_sc_hd__buf_2
XFILLER_204_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_82_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_82_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19279_ _19837_/A _20149_/B _19278_/X VGND VGND VPWR VPWR _19280_/A sky130_fd_sc_hd__or3_4
XFILLER_175_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21310_ _15866_/X VGND VGND VPWR VPWR _21311_/A sky130_fd_sc_hd__buf_2
XFILLER_163_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22290_ _21719_/B VGND VGND VPWR VPWR _22291_/B sky130_fd_sc_hd__buf_2
XANTENNA__16516__A1_N _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21241_ _21273_/A _21241_/B VGND VGND VPWR VPWR _21244_/B sky130_fd_sc_hd__or2_4
XFILLER_190_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14226__A2_N _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21172_ _16864_/Y _21172_/B VGND VGND VPWR VPWR _21175_/B sky130_fd_sc_hd__or2_4
XFILLER_172_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20123_ _21418_/B _20118_/X _20122_/X _20118_/X VGND VGND VPWR VPWR _23510_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17128__A _17074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19416__B1 _19326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21873__A _16731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22566__A3 _22145_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20054_ _21477_/B _20051_/X _20010_/X _20051_/X VGND VGND VPWR VPWR _23534_/D sky130_fd_sc_hd__a2bb2o_4
X_24931_ _23678_/CLK _24931_/D HRESETn VGND VGND VPWR VPWR _13603_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_140_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24862_ _24476_/CLK _24862_/D HRESETn VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23813_ _23454_/CLK _19255_/X VGND VGND VPWR VPWR _23813_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24793_ _24825_/CLK _15915_/X HRESETn VGND VGND VPWR VPWR _21712_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23754_/CLK _23744_/D VGND VGND VPWR VPWR _18118_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _20956_/A VGND VGND VPWR VPWR _20956_/Y sky130_fd_sc_hd__inv_2
XPHY_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_31_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23644_/CLK _19657_/X VGND VGND VPWR VPWR _13251_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _20878_/X _20886_/X _16701_/A _20883_/X VGND VGND VPWR VPWR _20887_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _16432_/A _22589_/B VGND VGND VPWR VPWR _22629_/B sky130_fd_sc_hd__or2_4
X_25414_ _24867_/CLK _12726_/X HRESETn VGND VGND VPWR VPWR _25414_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25148__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11778__B1 _11776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25345_ _25368_/CLK _25345_/D HRESETn VGND VGND VPWR VPWR _12351_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21113__A _21064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22557_ _22557_/A _16382_/A VGND VGND VPWR VPWR _22561_/B sky130_fd_sc_hd__or2_4
XFILLER_166_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16207__A _23218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12310_ _12310_/A _12310_/B _12307_/X _12310_/D VGND VGND VPWR VPWR _12310_/X sky130_fd_sc_hd__or4_4
X_21508_ _21503_/X _21507_/X _18306_/X VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__o21a_4
X_13290_ _13451_/A VGND VGND VPWR VPWR _13290_/X sky130_fd_sc_hd__buf_2
X_25276_ _25276_/CLK _25276_/D HRESETn VGND VGND VPWR VPWR _25276_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12990__A2 _12875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22488_ _21430_/X VGND VGND VPWR VPWR _22488_/X sky130_fd_sc_hd__buf_2
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ _22159_/A VGND VGND VPWR VPWR _12241_/Y sky130_fd_sc_hd__inv_2
X_24227_ _24206_/CLK _24227_/D HRESETn VGND VGND VPWR VPWR _21514_/A sky130_fd_sc_hd__dfrtp_4
X_21439_ _22430_/A _21439_/B VGND VGND VPWR VPWR _21439_/Y sky130_fd_sc_hd__nand2_4
XFILLER_107_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _12170_/X _12172_/B VGND VGND VPWR VPWR _12172_/X sky130_fd_sc_hd__and2_4
X_24158_ _24160_/CLK _24158_/D HRESETn VGND VGND VPWR VPWR _24158_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23109_ _22771_/X _23107_/X _22702_/X _23108_/X VGND VGND VPWR VPWR _23110_/A sky130_fd_sc_hd__o22a_4
XFILLER_122_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22006__A2 _20356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16980_ _16973_/X _16980_/B _16980_/C _16979_/X VGND VGND VPWR VPWR _16980_/X sky130_fd_sc_hd__or4_4
X_24089_ _23980_/CLK _24089_/D HRESETn VGND VGND VPWR VPWR _24089_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21555__A1_N _17389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15931_ _15659_/B _15934_/B VGND VGND VPWR VPWR _15931_/X sky130_fd_sc_hd__or2_4
XFILLER_89_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17969__B1 _15686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16877__A _14791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15781__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18650_ _16601_/Y _18693_/A _16601_/Y _18693_/A VGND VGND VPWR VPWR _18650_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15862_ _21589_/B VGND VGND VPWR VPWR _22684_/B sky130_fd_sc_hd__buf_2
XFILLER_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17601_ _17566_/Y _17595_/B _17596_/B _17600_/X VGND VGND VPWR VPWR _17601_/X sky130_fd_sc_hd__a211o_4
X_14813_ _14812_/X VGND VGND VPWR VPWR _14815_/B sky130_fd_sc_hd__inv_2
X_18581_ _18556_/X _18572_/B _18581_/C VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__and3_4
X_15793_ _14386_/A _15792_/X VGND VGND VPWR VPWR _15793_/X sky130_fd_sc_hd__or2_4
XFILLER_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22714__B1 _15676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24680__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17532_ _25543_/Q _17531_/A _11796_/Y _17531_/Y VGND VGND VPWR VPWR _17532_/X sky130_fd_sc_hd__o22a_4
XFILLER_123_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14744_ _22060_/A _14717_/X _25073_/Q _14715_/X VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__o22a_4
X_11956_ _11934_/X VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__buf_2
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18394__B1 _24196_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17463_ _17464_/A VGND VGND VPWR VPWR _17463_/X sky130_fd_sc_hd__buf_2
XFILLER_199_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11887_ _11887_/A _11887_/B VGND VGND VPWR VPWR _11887_/Y sky130_fd_sc_hd__nand2_4
X_14675_ _19054_/A _14668_/X _14674_/X VGND VGND VPWR VPWR _25079_/D sky130_fd_sc_hd__a21oi_4
XANTENNA__18605__A1_N _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19202_ _23831_/Q VGND VGND VPWR VPWR _19202_/Y sky130_fd_sc_hd__inv_2
X_16414_ HWDATA[19] VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__buf_2
X_13626_ _13626_/A VGND VGND VPWR VPWR _13628_/A sky130_fd_sc_hd__inv_2
XANTENNA__23222__B _23313_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17394_ _17353_/A _17391_/B _17393_/X VGND VGND VPWR VPWR _24346_/D sky130_fd_sc_hd__and3_4
XFILLER_158_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19133_ _23855_/Q VGND VGND VPWR VPWR _19133_/Y sky130_fd_sc_hd__inv_2
X_16345_ _24628_/Q VGND VGND VPWR VPWR _16345_/Y sky130_fd_sc_hd__inv_2
X_13557_ _25094_/Q VGND VGND VPWR VPWR _14607_/A sky130_fd_sc_hd__inv_2
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12508_ _12232_/Y _12514_/B VGND VGND VPWR VPWR _12508_/X sky130_fd_sc_hd__or2_4
X_19064_ _19063_/Y _19061_/X _18969_/X _19061_/X VGND VGND VPWR VPWR _23881_/D sky130_fd_sc_hd__a2bb2o_4
X_13488_ _25328_/Q VGND VGND VPWR VPWR _13488_/Y sky130_fd_sc_hd__inv_2
X_16276_ _14479_/A VGND VGND VPWR VPWR _16276_/X sky130_fd_sc_hd__buf_2
X_18015_ _18130_/A _18012_/X _18015_/C VGND VGND VPWR VPWR _18016_/C sky130_fd_sc_hd__and3_4
X_12439_ _12439_/A _12439_/B _12292_/X _12391_/X VGND VGND VPWR VPWR _12440_/C sky130_fd_sc_hd__or4_4
X_15227_ _15227_/A VGND VGND VPWR VPWR _25033_/D sky130_fd_sc_hd__inv_2
XFILLER_173_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12194__B1 _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21453__B1 _12353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15158_ _15158_/A VGND VGND VPWR VPWR _15158_/Y sky130_fd_sc_hd__inv_2
X_14109_ _25221_/Q _14109_/B _14124_/A VGND VGND VPWR VPWR _14110_/B sky130_fd_sc_hd__or3_4
X_15089_ _25006_/Q VGND VGND VPWR VPWR _15303_/A sky130_fd_sc_hd__inv_2
X_19966_ _19965_/X VGND VGND VPWR VPWR _19979_/A sky130_fd_sc_hd__inv_2
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22789__A _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18917_ _18916_/Y VGND VGND VPWR VPWR _18917_/X sky130_fd_sc_hd__buf_2
XANTENNA__21693__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19897_ _19897_/A VGND VGND VPWR VPWR _21474_/B sky130_fd_sc_hd__inv_2
XFILLER_122_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24768__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _16472_/A _24161_/Q _16472_/Y _18678_/Y VGND VGND VPWR VPWR _18850_/C sky130_fd_sc_hd__o22a_4
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16632__B1 _16375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18779_ _18710_/A _18700_/A VGND VGND VPWR VPWR _18779_/X sky130_fd_sc_hd__or2_4
XFILLER_227_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20810_ _13127_/B _20809_/A VGND VGND VPWR VPWR _20810_/X sky130_fd_sc_hd__or2_4
X_21790_ _21644_/A _21790_/B VGND VGND VPWR VPWR _21790_/X sky130_fd_sc_hd__or2_4
XANTENNA__13642__C _13636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17188__B2 _17294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16440__A1_N _15108_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20741_ _13139_/A _13138_/X _20740_/Y VGND VGND VPWR VPWR _20741_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23460_ _23459_/CLK _23460_/D VGND VGND VPWR VPWR _20255_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20672_ _20672_/A _17413_/A VGND VGND VPWR VPWR _20675_/B sky130_fd_sc_hd__or2_4
XFILLER_189_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22029__A _22029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22411_ _22541_/A VGND VGND VPWR VPWR _22411_/X sky130_fd_sc_hd__buf_2
X_23391_ _23913_/CLK _20431_/X VGND VGND VPWR VPWR _13316_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_176_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25556__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15539__A2_N _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25130_ _25125_/CLK _14473_/X HRESETn VGND VGND VPWR VPWR _25130_/Q sky130_fd_sc_hd__dfrtp_4
X_22342_ _21350_/Y _22327_/X _22329_/X _22333_/Y _22341_/X VGND VGND VPWR VPWR _22401_/C
+ sky130_fd_sc_hd__a2111o_4
XFILLER_149_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25061_ _23385_/CLK _14830_/X HRESETn VGND VGND VPWR VPWR _25061_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15866__A _21173_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22273_ _18301_/A _22269_/X _22272_/X VGND VGND VPWR VPWR _22273_/X sky130_fd_sc_hd__or3_4
XFILLER_164_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12185__B1 _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24012_ _24012_/CLK _20531_/X HRESETn VGND VGND VPWR VPWR _20530_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_26_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _24937_/CLK sky130_fd_sc_hd__clkbuf_1
X_21224_ _21224_/A VGND VGND VPWR VPWR _21224_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_89_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _24856_/CLK sky130_fd_sc_hd__clkbuf_1
X_21155_ _21155_/A _21154_/X VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__and2_4
XFILLER_160_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23197__B1 _24852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20106_ _20104_/Y _20101_/X _20105_/X _20101_/X VGND VGND VPWR VPWR _20106_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21086_ _21172_/B VGND VGND VPWR VPWR _21231_/A sky130_fd_sc_hd__buf_2
X_20037_ _17717_/X _18293_/X _18290_/A _19986_/X VGND VGND VPWR VPWR _20038_/A sky130_fd_sc_hd__or4_4
X_24914_ _24915_/CLK _24914_/D HRESETn VGND VGND VPWR VPWR _24914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24845_ _24849_/CLK _24845_/D HRESETn VGND VGND VPWR VPWR _24845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11807_/Y _11804_/X _11809_/X _11804_/X VGND VGND VPWR VPWR _25540_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A VGND VGND VPWR VPWR _12790_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _21282_/X _21986_/X _21987_/X _23358_/A _21654_/X VGND VGND VPWR VPWR _21989_/B
+ sky130_fd_sc_hd__a32o_4
X_24776_ _24803_/CLK _24776_/D HRESETn VGND VGND VPWR VPWR _23049_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_15_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _15661_/C VGND VGND VPWR VPWR _21045_/A sky130_fd_sc_hd__buf_2
XFILLER_82_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20939_ _20939_/A VGND VGND VPWR VPWR _20939_/Y sky130_fd_sc_hd__inv_2
X_23727_ _23717_/CLK _19497_/X VGND VGND VPWR VPWR _23727_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16926__B2 _16925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11672_/A VGND VGND VPWR VPWR _11672_/Y sky130_fd_sc_hd__inv_2
X_14460_ _14191_/Y _14457_/X _14409_/X _14446_/A VGND VGND VPWR VPWR _25135_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _23642_/CLK _23658_/D VGND VGND VPWR VPWR _13288_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13411_/A _13411_/B VGND VGND VPWR VPWR _13411_/X sky130_fd_sc_hd__or2_4
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _14390_/B _14389_/X _14392_/A VGND VGND VPWR VPWR _14391_/X sky130_fd_sc_hd__a21o_4
X_22609_ _22494_/X _22608_/X _21303_/A _24836_/Q _22569_/X VGND VGND VPWR VPWR _22609_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23589_ _23565_/CLK _23589_/D VGND VGND VPWR VPWR _23589_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13342_ _13187_/X _13331_/X _13341_/X VGND VGND VPWR VPWR _13342_/X sky130_fd_sc_hd__and3_4
X_16130_ _22883_/A VGND VGND VPWR VPWR _16130_/Y sky130_fd_sc_hd__inv_2
X_25328_ _24112_/CLK _25328_/D HRESETn VGND VGND VPWR VPWR _25328_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20682__A _20686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13273_ _13412_/A _13270_/X _13273_/C VGND VGND VPWR VPWR _13277_/B sky130_fd_sc_hd__and3_4
X_16061_ _16044_/A VGND VGND VPWR VPWR _16061_/X sky130_fd_sc_hd__buf_2
X_25259_ _25204_/CLK _25259_/D HRESETn VGND VGND VPWR VPWR _13862_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12224_ _25457_/Q _22910_/A _12222_/Y _12223_/Y VGND VGND VPWR VPWR _12224_/X sky130_fd_sc_hd__o22a_4
X_15012_ _15012_/A VGND VGND VPWR VPWR _15012_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19820_ _19819_/Y _19816_/X _19769_/X _19816_/X VGND VGND VPWR VPWR _23619_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13296__A _13320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12155_ _12140_/A _20982_/A _12140_/Y _12154_/X VGND VGND VPWR VPWR _12166_/A sky130_fd_sc_hd__a211o_4
XANTENNA__17991__A _18097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11809__A _16238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16862__B1 _16861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19751_ _19750_/Y _19748_/X _19728_/X _19748_/X VGND VGND VPWR VPWR _19751_/X sky130_fd_sc_hd__a2bb2o_4
X_12086_ _12085_/Y _12083_/X _11847_/X _12083_/X VGND VGND VPWR VPWR _12086_/X sky130_fd_sc_hd__a2bb2o_4
X_16963_ _16962_/X VGND VGND VPWR VPWR _16963_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24861__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18702_ _18702_/A _18701_/X VGND VGND VPWR VPWR _18702_/X sky130_fd_sc_hd__or2_4
X_15914_ _15714_/X _15902_/X _15775_/X _24794_/Q _15871_/X VGND VGND VPWR VPWR _15914_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19682_ _19675_/Y VGND VGND VPWR VPWR _19682_/X sky130_fd_sc_hd__buf_2
X_16894_ _16887_/X VGND VGND VPWR VPWR _16894_/X sky130_fd_sc_hd__buf_2
XFILLER_65_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16614__B1 _16613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _24150_/Q VGND VGND VPWR VPWR _18698_/C sky130_fd_sc_hd__inv_2
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15845_ _15833_/X _15844_/X _15775_/X _24829_/Q _15802_/A VGND VGND VPWR VPWR _24829_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18564_ _18564_/A VGND VGND VPWR VPWR _24175_/D sky130_fd_sc_hd__inv_2
XANTENNA__19711__A _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15776_ _15758_/X _15774_/X _15775_/X _24864_/Q _15719_/X VGND VGND VPWR VPWR _15776_/X
+ sky130_fd_sc_hd__a32o_4
X_12988_ _12988_/A _12988_/B _12988_/C VGND VGND VPWR VPWR _25373_/D sky130_fd_sc_hd__and3_4
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22163__A1 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12100__B1 _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22163__B2 _22947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17515_ _17515_/A _17510_/X _17513_/X _17515_/D VGND VGND VPWR VPWR _17515_/X sky130_fd_sc_hd__or4_4
X_14727_ _14725_/X _14726_/X _14725_/X _14726_/X VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__a2bb2o_4
X_11939_ _19626_/A VGND VGND VPWR VPWR _11939_/X sky130_fd_sc_hd__buf_2
X_18495_ _18489_/A _18488_/X _18490_/B _18494_/X VGND VGND VPWR VPWR _18496_/A sky130_fd_sc_hd__a211o_4
XFILLER_221_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _17445_/Y _17441_/X _16729_/X _17426_/A VGND VGND VPWR VPWR _24331_/D sky130_fd_sc_hd__a2bb2o_4
X_14658_ _25080_/Q VGND VGND VPWR VPWR _17985_/A sky130_fd_sc_hd__inv_2
XFILLER_21_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13609_ _14668_/A VGND VGND VPWR VPWR _19054_/D sky130_fd_sc_hd__inv_2
X_17377_ _17198_/X _17375_/X _17376_/Y VGND VGND VPWR VPWR _17377_/X sky130_fd_sc_hd__o21a_4
X_14589_ _14588_/X VGND VGND VPWR VPWR _14590_/B sky130_fd_sc_hd__inv_2
X_19116_ _23861_/Q VGND VGND VPWR VPWR _19116_/Y sky130_fd_sc_hd__inv_2
X_16328_ _16327_/Y _16325_/X _15970_/X _16325_/X VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_185_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11710__C _11889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17185__A1_N _16348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19047_ HWDATA[1] VGND VGND VPWR VPWR _19048_/A sky130_fd_sc_hd__buf_2
XFILLER_146_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16259_ _24660_/Q VGND VGND VPWR VPWR _16259_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_242_0_HCLK clkbuf_8_242_0_HCLK/A VGND VGND VPWR VPWR _25212_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20229__B2 _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11719__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19949_ _22264_/B _19946_/X _19629_/X _19946_/X VGND VGND VPWR VPWR _23571_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21729__A1 _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22960_ _22836_/A _22960_/B _22960_/C VGND VGND VPWR VPWR _22979_/B sky130_fd_sc_hd__and3_4
XANTENNA__24531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16605__B1 _16252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21911_ _22373_/A _21909_/X _21911_/C VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__and3_4
X_22891_ _15601_/Y _22891_/B VGND VGND VPWR VPWR _22891_/X sky130_fd_sc_hd__and2_4
XFILLER_215_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21842_ _24051_/Q VGND VGND VPWR VPWR _21842_/Y sky130_fd_sc_hd__inv_2
X_24630_ _24629_/CLK _24630_/D HRESETn VGND VGND VPWR VPWR _24630_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21870__B _21855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24561_ _24528_/CLK _16526_/X HRESETn VGND VGND VPWR VPWR _24561_/Q sky130_fd_sc_hd__dfrtp_4
X_21773_ _14761_/A _21773_/B VGND VGND VPWR VPWR _21773_/X sky130_fd_sc_hd__or2_4
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16908__B2 _24289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20724_/A VGND VGND VPWR VPWR _20724_/X sky130_fd_sc_hd__buf_2
X_23512_ _23513_/CLK _23512_/D VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24492_ _24493_/CLK _16710_/X HRESETn VGND VGND VPWR VPWR _16708_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _23555_/CLK _23443_/D VGND VGND VPWR VPWR _20300_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20655_ _20654_/X VGND VGND VPWR VPWR _20655_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_52_0_HCLK clkbuf_5_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23374_ _23361_/X VGND VGND VPWR VPWR IRQ[18] sky130_fd_sc_hd__buf_2
X_20586_ _14437_/Y _20574_/X _20565_/X _20585_/X VGND VGND VPWR VPWR _20587_/A sky130_fd_sc_hd__a211o_4
X_22325_ _22324_/Y _21353_/X _14414_/Y _21356_/X VGND VGND VPWR VPWR _22326_/A sky130_fd_sc_hd__o22a_4
X_25113_ _23970_/CLK _14529_/X HRESETn VGND VGND VPWR VPWR _25113_/Q sky130_fd_sc_hd__dfrtp_4
X_25044_ _25043_/CLK _25044_/D HRESETn VGND VGND VPWR VPWR _14897_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_219_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22256_ _22264_/A _22256_/B VGND VGND VPWR VPWR _22256_/X sky130_fd_sc_hd__or2_4
XANTENNA__13828__B _13782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21207_ _21207_/A _20381_/Y VGND VGND VPWR VPWR _21209_/B sky130_fd_sc_hd__or2_4
X_22187_ _12118_/Y _12107_/A _18381_/Y _12080_/A VGND VGND VPWR VPWR _22187_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23963__D scl_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24619__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16844__B1 _15759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21138_ _14408_/Y _21861_/A _14481_/Y _21373_/A VGND VGND VPWR VPWR _21138_/X sky130_fd_sc_hd__o22a_4
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17316__A _17257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13960_ _13952_/D VGND VGND VPWR VPWR _13960_/Y sky130_fd_sc_hd__inv_2
X_21069_ _21069_/A _21069_/B VGND VGND VPWR VPWR _21069_/X sky130_fd_sc_hd__or2_4
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23037__B _22968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _22678_/A _12941_/A _12609_/X _12856_/X VGND VGND VPWR VPWR _12911_/X sky130_fd_sc_hd__or4_4
XFILLER_207_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13891_ _21160_/A _13869_/X _23444_/Q _13864_/X VGND VGND VPWR VPWR _13891_/X sky130_fd_sc_hd__o22a_4
XFILLER_246_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15630_ _15628_/Y _15626_/X _15629_/X _15626_/X VGND VGND VPWR VPWR _15630_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12842_ _12842_/A VGND VGND VPWR VPWR _12969_/A sky130_fd_sc_hd__inv_2
X_24828_ _24825_/CLK _15846_/X HRESETn VGND VGND VPWR VPWR _24828_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23053__A _23053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15561_ _15560_/X VGND VGND VPWR VPWR _15561_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12773_ _12773_/A VGND VGND VPWR VPWR _12773_/Y sky130_fd_sc_hd__inv_2
X_24759_ _24759_/CLK _15989_/X HRESETn VGND VGND VPWR VPWR _22285_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17231_/Y _17265_/X _17355_/B VGND VGND VPWR VPWR _17300_/X sky130_fd_sc_hd__or3_4
XANTENNA__17021__B1 _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _25117_/Q _14517_/A VGND VGND VPWR VPWR _14512_/Y sky130_fd_sc_hd__nor2_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11724_ _11724_/A VGND VGND VPWR VPWR _15791_/C sky130_fd_sc_hd__buf_2
X_18280_ _13793_/D _20408_/A _13481_/A _24225_/Q _18279_/X VGND VGND VPWR VPWR _24225_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15492_/A VGND VGND VPWR VPWR _15493_/B sky130_fd_sc_hd__inv_2
XFILLER_70_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A VGND VGND VPWR VPWR _17231_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443_ _14443_/A VGND VGND VPWR VPWR _22334_/B sky130_fd_sc_hd__buf_2
XANTENNA__17986__A _18008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22448__A2 _22425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _17162_/A VGND VGND VPWR VPWR _17162_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25204__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14374_ _14364_/X _14373_/X _12090_/A _14369_/X VGND VGND VPWR VPWR _14374_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _24711_/Q VGND VGND VPWR VPWR _16113_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21301__A _21300_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13325_ _13286_/X _13325_/B VGND VGND VPWR VPWR _13325_/X sky130_fd_sc_hd__or2_4
XFILLER_116_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15335__B1 _15324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17093_ _17093_/A VGND VGND VPWR VPWR _17094_/B sky130_fd_sc_hd__inv_2
XFILLER_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16044_ _16044_/A VGND VGND VPWR VPWR _16044_/X sky130_fd_sc_hd__buf_2
X_13256_ _13428_/A _19722_/A VGND VGND VPWR VPWR _13256_/X sky130_fd_sc_hd__or2_4
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _12198_/X _12207_/B _12204_/X _12206_/X VGND VGND VPWR VPWR _12207_/X sky130_fd_sc_hd__or4_4
X_13187_ _13186_/Y VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_72_0_HCLK clkbuf_8_73_0_HCLK/A VGND VGND VPWR VPWR _24712_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16835__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _12138_/A VGND VGND VPWR VPWR _12138_/Y sky130_fd_sc_hd__inv_2
X_19803_ _19803_/A VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__buf_2
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17995_ _18178_/A _17995_/B VGND VGND VPWR VPWR _17995_/X sky130_fd_sc_hd__or2_4
XFILLER_215_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12069_ _13484_/C _12081_/B _13542_/C _12068_/X VGND VGND VPWR VPWR _12070_/A sky130_fd_sc_hd__or4_4
X_16946_ _16942_/X _16943_/X _16944_/X _16945_/X VGND VGND VPWR VPWR _16946_/X sky130_fd_sc_hd__or4_4
X_19734_ _11865_/X VGND VGND VPWR VPWR _19734_/X sky130_fd_sc_hd__buf_2
XFILLER_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19665_ _19664_/Y _19660_/X _19612_/X _19660_/X VGND VGND VPWR VPWR _23672_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16877_ _14791_/X VGND VGND VPWR VPWR _16877_/X sky130_fd_sc_hd__buf_2
X_18616_ _16606_/A _18794_/C _16566_/Y _24157_/Q VGND VGND VPWR VPWR _18616_/X sky130_fd_sc_hd__a2bb2o_4
X_15828_ _15844_/A VGND VGND VPWR VPWR _15828_/X sky130_fd_sc_hd__buf_2
X_19596_ _21380_/A VGND VGND VPWR VPWR _21382_/C sky130_fd_sc_hd__inv_2
XANTENNA__23333__B1 _25404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18547_ _18540_/B _18550_/B VGND VGND VPWR VPWR _18548_/C sky130_fd_sc_hd__nand2_4
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15759_ HWDATA[12] VGND VGND VPWR VPWR _15759_/X sky130_fd_sc_hd__buf_2
XFILLER_178_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18478_ _24174_/Q VGND VGND VPWR VPWR _18479_/C sky130_fd_sc_hd__inv_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _17429_/A VGND VGND VPWR VPWR _17429_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20440_ _14389_/B VGND VGND VPWR VPWR _20463_/C sky130_fd_sc_hd__inv_2
XFILLER_158_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20371_ _20369_/Y _20365_/X _19632_/A _20370_/X VGND VGND VPWR VPWR _20371_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22110_ _16620_/A _22299_/B _22108_/X _22109_/X VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__a211o_4
XFILLER_146_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23090_ _17195_/A _21034_/X VGND VGND VPWR VPWR _23093_/B sky130_fd_sc_hd__or2_4
XFILLER_161_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24783__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22041_ _21682_/A _22041_/B VGND VGND VPWR VPWR _22041_/X sky130_fd_sc_hd__or2_4
XANTENNA__17618__A2 _17610_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22611__A2 _22610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24712__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16826__B1 HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23021__C1 _23020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23992_ _23991_/CLK _20650_/Y HRESETn VGND VGND VPWR VPWR _17401_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16040__A _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22943_ _24539_/Q _22940_/X _22941_/X _22942_/X VGND VGND VPWR VPWR _22944_/C sky130_fd_sc_hd__a211o_4
XFILLER_29_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22874_ _22487_/A _22873_/X VGND VGND VPWR VPWR _22874_/X sky130_fd_sc_hd__and2_4
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24613_ _24613_/CLK _24613_/D HRESETn VGND VGND VPWR VPWR _24613_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21825_ _21687_/A _21825_/B VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__or2_4
XFILLER_231_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21756_ _16720_/Y _22575_/A VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__and2_4
X_24544_ _24542_/CLK _24544_/D HRESETn VGND VGND VPWR VPWR _16571_/A sky130_fd_sc_hd__dfrtp_4
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21886__B1 _11853_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _20706_/X VGND VGND VPWR VPWR _20707_/Y sky130_fd_sc_hd__inv_2
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21687_ _21687_/A _19916_/Y VGND VGND VPWR VPWR _21689_/B sky130_fd_sc_hd__or2_4
X_24475_ _24473_/CLK _24475_/D HRESETn VGND VGND VPWR VPWR _15051_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20638_ _17399_/A _17399_/B VGND VGND VPWR VPWR _20639_/B sky130_fd_sc_hd__nand2_4
X_23426_ _23400_/CLK _23426_/D VGND VGND VPWR VPWR _22275_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21121__A _21121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23357_ _18273_/Y _21834_/A _17490_/Y _21514_/A VGND VGND VPWR VPWR _23357_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20569_ _20569_/A VGND VGND VPWR VPWR _23952_/D sky130_fd_sc_hd__inv_2
XFILLER_153_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13110_ _13091_/B VGND VGND VPWR VPWR _13111_/B sky130_fd_sc_hd__inv_2
X_22308_ _22307_/Y _22296_/X _24021_/Q _21296_/X VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__a2bb2o_4
X_14090_ _14082_/A VGND VGND VPWR VPWR _14090_/X sky130_fd_sc_hd__buf_2
X_23288_ _23113_/X _23287_/X _23159_/X _24855_/Q _23115_/X VGND VGND VPWR VPWR _23288_/X
+ sky130_fd_sc_hd__a32o_4
X_13041_ _12308_/Y _13044_/B _13040_/X VGND VGND VPWR VPWR _13041_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_124_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22239_ _19554_/A _22013_/Y _22524_/B _22238_/X VGND VGND VPWR VPWR _22240_/A sky130_fd_sc_hd__a211o_4
X_25027_ _25023_/CLK _15246_/Y HRESETn VGND VGND VPWR VPWR _14958_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22602__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16817__B1 _15732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_59_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23048__A _23025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16800_ _16799_/Y _16738_/X _16726_/X _16738_/X VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17780_ _16962_/X _17609_/B VGND VGND VPWR VPWR _17780_/X sky130_fd_sc_hd__and2_4
X_14992_ _14985_/X _14987_/X _14988_/X _14991_/X VGND VGND VPWR VPWR _14992_/X sky130_fd_sc_hd__or4_4
XFILLER_247_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16731_ _16379_/A VGND VGND VPWR VPWR _16731_/Y sky130_fd_sc_hd__inv_2
X_13943_ _13942_/X _13934_/X _13899_/C _13948_/C VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__or4_4
XFILLER_219_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19450_ _18150_/B VGND VGND VPWR VPWR _19450_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16662_ _16662_/A VGND VGND VPWR VPWR _16662_/Y sky130_fd_sc_hd__inv_2
X_13874_ _13861_/X _13873_/X VGND VGND VPWR VPWR _13874_/X sky130_fd_sc_hd__or2_4
X_18401_ _16263_/A _18400_/Y _16207_/Y _24190_/Q VGND VGND VPWR VPWR _18401_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23315__B1 _22815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15613_ _24911_/Q VGND VGND VPWR VPWR _15613_/Y sky130_fd_sc_hd__inv_2
X_12825_ _25395_/Q VGND VGND VPWR VPWR _12825_/Y sky130_fd_sc_hd__inv_2
X_19381_ _18142_/B VGND VGND VPWR VPWR _19381_/Y sky130_fd_sc_hd__inv_2
X_16593_ _16590_/Y _16592_/X _16334_/X _16592_/X VGND VGND VPWR VPWR _24536_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12606__B2 _24863_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18332_ _18332_/A VGND VGND VPWR VPWR _19075_/B sky130_fd_sc_hd__buf_2
XFILLER_188_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11822__A _16248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15544_ _15544_/A VGND VGND VPWR VPWR _15544_/X sky130_fd_sc_hd__buf_2
X_12756_ _12888_/A VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__inv_2
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11705_/A _24244_/Q _11705_/Y _11706_/Y VGND VGND VPWR VPWR _11708_/D sky130_fd_sc_hd__o22a_4
X_18263_ _13828_/D _18262_/X _15993_/X _24234_/Q _18248_/A VGND VGND VPWR VPWR _24234_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15474_/Y _15472_/X _14423_/X _15472_/X VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12687_ _12618_/A _12691_/B _12686_/Y VGND VGND VPWR VPWR _12687_/X sky130_fd_sc_hd__o21a_4
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _24347_/Q VGND VGND VPWR VPWR _17214_/Y sky130_fd_sc_hd__inv_2
X_14426_ HWDATA[5] VGND VGND VPWR VPWR _14427_/A sky130_fd_sc_hd__buf_2
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18194_ _18063_/A _18194_/B _18194_/C VGND VGND VPWR VPWR _18195_/C sky130_fd_sc_hd__and3_4
XANTENNA__23094__A2 _21890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16854__A1_N _14899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17050_/C _17144_/X _17065_/X VGND VGND VPWR VPWR _17145_/Y sky130_fd_sc_hd__a21oi_4
X_14357_ _14352_/X VGND VGND VPWR VPWR _14360_/A sky130_fd_sc_hd__inv_2
X_13308_ _13411_/A _23857_/Q VGND VGND VPWR VPWR _13309_/C sky130_fd_sc_hd__or2_4
XANTENNA__21966__A _22274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17076_ _17393_/B VGND VGND VPWR VPWR _17076_/X sky130_fd_sc_hd__buf_2
XFILLER_116_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14288_ _15465_/A VGND VGND VPWR VPWR _15446_/A sky130_fd_sc_hd__buf_2
X_16027_ _16026_/Y _16024_/X _11780_/X _16024_/X VGND VGND VPWR VPWR _16027_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13239_ _13391_/A _13239_/B _13239_/C VGND VGND VPWR VPWR _13240_/C sky130_fd_sc_hd__or3_4
XFILLER_226_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17978_ _17985_/A VGND VGND VPWR VPWR _17979_/A sky130_fd_sc_hd__buf_2
XFILLER_111_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16929_ _16929_/A VGND VGND VPWR VPWR _16929_/Y sky130_fd_sc_hd__inv_2
X_19717_ _13173_/B VGND VGND VPWR VPWR _19717_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16795__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19648_ _19648_/A VGND VGND VPWR VPWR _21195_/B sky130_fd_sc_hd__inv_2
XANTENNA__22109__A1 _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19579_ _23698_/Q VGND VGND VPWR VPWR _22041_/B sky130_fd_sc_hd__inv_2
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21610_ _21564_/Y _21610_/B _21610_/C _21609_/X VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__or4_4
XANTENNA__18218__C _18217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22590_ _24462_/Q _22543_/X _22544_/X VGND VGND VPWR VPWR _22590_/X sky130_fd_sc_hd__o21a_4
XFILLER_240_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21541_ _15792_/X VGND VGND VPWR VPWR _21542_/A sky130_fd_sc_hd__buf_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18515__A _18515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21883__A3 _22954_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24260_ _23494_/CLK _24260_/D HRESETn VGND VGND VPWR VPWR _22003_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21472_ _21472_/A VGND VGND VPWR VPWR _21482_/A sky130_fd_sc_hd__buf_2
XANTENNA__19289__B2 _19286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23211_ _23209_/X _23210_/X _22150_/A VGND VGND VPWR VPWR _23211_/X sky130_fd_sc_hd__or3_4
XANTENNA__24101__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20423_ _20430_/A VGND VGND VPWR VPWR _20423_/X sky130_fd_sc_hd__buf_2
X_24191_ _24194_/CLK _18507_/Y HRESETn VGND VGND VPWR VPWR _24191_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22293__B1 _22836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23142_ _23136_/X _23142_/B VGND VGND VPWR VPWR _23142_/Y sky130_fd_sc_hd__nor2_4
X_20354_ _23423_/Q VGND VGND VPWR VPWR _21995_/B sky130_fd_sc_hd__buf_2
XFILLER_162_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23073_ _20797_/Y _23006_/X _20936_/Y _21229_/X VGND VGND VPWR VPWR _23073_/X sky130_fd_sc_hd__o22a_4
X_20285_ _22085_/B _20279_/X _16874_/X _20284_/X VGND VGND VPWR VPWR _23450_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22024_ _22032_/A _20307_/Y VGND VGND VPWR VPWR _22025_/C sky130_fd_sc_hd__or2_4
XFILLER_103_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13394__A _13282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20359__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23975_ _23385_/CLK _25189_/Q HRESETn VGND VGND VPWR VPWR _22338_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22899__A2 _21085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22926_ _22437_/X VGND VGND VPWR VPWR _22926_/X sky130_fd_sc_hd__buf_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18972__B1 _16796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22857_ _22837_/X _22841_/Y _22848_/Y _22856_/X VGND VGND VPWR VPWR _22870_/C sky130_fd_sc_hd__a211o_4
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12610_ _12609_/X VGND VGND VPWR VPWR _12638_/B sky130_fd_sc_hd__buf_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12352__A2_N _12350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15114__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21808_ _21808_/A _21806_/X _21807_/X VGND VGND VPWR VPWR _21808_/X sky130_fd_sc_hd__and3_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590_ _13840_/A _14601_/A _13589_/Y _25098_/Q VGND VGND VPWR VPWR _13590_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22788_ _22721_/B VGND VGND VPWR VPWR _22788_/X sky130_fd_sc_hd__buf_2
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12541_ _12541_/A VGND VGND VPWR VPWR _12618_/A sky130_fd_sc_hd__inv_2
X_24527_ _24556_/CLK _16616_/X HRESETn VGND VGND VPWR VPWR _16615_/A sky130_fd_sc_hd__dfrtp_4
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21739_ _21732_/Y _21733_/Y _21739_/C _21739_/D VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__or4_4
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15260_ _15271_/A _15268_/A _15260_/C _15259_/X VGND VGND VPWR VPWR _15260_/X sky130_fd_sc_hd__or4_4
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12472_ _12439_/A _12469_/X VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__or2_4
X_24458_ _24425_/CLK _16786_/X HRESETn VGND VGND VPWR VPWR _24458_/Q sky130_fd_sc_hd__dfrtp_4
X_14211_ _20504_/A _14208_/X _13844_/X _14210_/X VGND VGND VPWR VPWR _14211_/X sky130_fd_sc_hd__a2bb2o_4
X_23409_ _23441_/CLK _23409_/D VGND VGND VPWR VPWR _20390_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_22_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_44_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15191_ _15182_/B _15181_/X _15183_/X _15188_/B VGND VGND VPWR VPWR _15191_/X sky130_fd_sc_hd__a211o_4
X_24389_ _24383_/CLK _17146_/X HRESETn VGND VGND VPWR VPWR _24389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24634__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14142_ _25228_/Q _14126_/X _14121_/Y _14128_/B VGND VGND VPWR VPWR _14142_/X sky130_fd_sc_hd__o22a_4
XFILLER_153_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14073_ _14073_/A VGND VGND VPWR VPWR _14082_/A sky130_fd_sc_hd__buf_2
X_18950_ _18949_/Y _18945_/X _16796_/X _18945_/X VGND VGND VPWR VPWR _23920_/D sky130_fd_sc_hd__a2bb2o_4
X_13024_ _13024_/A _13022_/A VGND VGND VPWR VPWR _13025_/C sky130_fd_sc_hd__or2_4
X_17901_ _17899_/A VGND VGND VPWR VPWR _17901_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18881_ _18881_/A _20571_/A VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__or2_4
XFILLER_239_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17832_ _17832_/A _17832_/B VGND VGND VPWR VPWR _17832_/X sky130_fd_sc_hd__or2_4
XANTENNA__11817__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17763_ _24275_/Q VGND VGND VPWR VPWR _17763_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14975_ _25017_/Q VGND VGND VPWR VPWR _15258_/A sky130_fd_sc_hd__inv_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_146_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _23647_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16714_ _16713_/Y _16709_/X _16534_/X _16709_/X VGND VGND VPWR VPWR _24490_/D sky130_fd_sc_hd__a2bb2o_4
X_19502_ _21190_/B _19496_/X _19501_/X _19483_/Y VGND VGND VPWR VPWR _23725_/D sky130_fd_sc_hd__a2bb2o_4
X_13926_ _13903_/Y _13921_/X _14260_/A VGND VGND VPWR VPWR _14254_/A sky130_fd_sc_hd__a21o_4
XFILLER_207_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17694_ _17538_/A _17693_/Y VGND VGND VPWR VPWR _17695_/B sky130_fd_sc_hd__or2_4
XANTENNA__23225__B _23222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19433_ _18213_/B VGND VGND VPWR VPWR _19433_/Y sky130_fd_sc_hd__inv_2
X_16645_ _16640_/A _16643_/X _16641_/Y _16644_/Y VGND VGND VPWR VPWR _16646_/A sky130_fd_sc_hd__a211o_4
X_13857_ _13857_/A VGND VGND VPWR VPWR _13857_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12648__A _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12808_ _12807_/Y VGND VGND VPWR VPWR _12941_/A sky130_fd_sc_hd__buf_2
X_19364_ _18224_/B VGND VGND VPWR VPWR _19364_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16576_ _16576_/A VGND VGND VPWR VPWR _16576_/Y sky130_fd_sc_hd__inv_2
X_13788_ _19595_/A _14228_/A VGND VGND VPWR VPWR _13789_/A sky130_fd_sc_hd__or2_4
X_18315_ _18314_/X VGND VGND VPWR VPWR _22271_/A sky130_fd_sc_hd__buf_2
X_15527_ _15524_/Y _15520_/X HADDR[12] _15526_/X VGND VGND VPWR VPWR _15527_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15529__B1 HADDR[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12739_ _12740_/A _12740_/B VGND VGND VPWR VPWR _12739_/Y sky130_fd_sc_hd__nand2_4
X_19295_ _23798_/Q VGND VGND VPWR VPWR _19295_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18246_ _20405_/A VGND VGND VPWR VPWR _20408_/A sky130_fd_sc_hd__inv_2
X_15458_ _15446_/A VGND VGND VPWR VPWR _15458_/X sky130_fd_sc_hd__buf_2
XANTENNA__21078__A1 _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14409_ _16729_/A VGND VGND VPWR VPWR _14409_/X sky130_fd_sc_hd__buf_2
X_18177_ _18039_/A _18177_/B VGND VGND VPWR VPWR _18177_/X sky130_fd_sc_hd__or2_4
XFILLER_117_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _15137_/Y _15389_/B VGND VGND VPWR VPWR _15390_/A sky130_fd_sc_hd__or2_4
XANTENNA__19140__B1 _19139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17128_ _17074_/A _17055_/C VGND VGND VPWR VPWR _17129_/B sky130_fd_sc_hd__or2_4
XFILLER_144_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21696__A _21815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17059_ _17074_/A _17072_/A _17034_/X _17068_/B VGND VGND VPWR VPWR _17059_/X sky130_fd_sc_hd__or4_4
XFILLER_116_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20070_ _21788_/B _20065_/X _19803_/X _20065_/X VGND VGND VPWR VPWR _23528_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_42_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22958__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20972_ _12010_/A _20972_/B VGND VGND VPWR VPWR _24104_/D sky130_fd_sc_hd__and2_4
X_23760_ _23768_/CLK _19403_/X VGND VGND VPWR VPWR _18111_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_226_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22711_ _22711_/A VGND VGND VPWR VPWR _22737_/B sky130_fd_sc_hd__inv_2
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23691_ _23690_/CLK _23691_/D VGND VGND VPWR VPWR _21981_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25430_ _25433_/CLK _25430_/D HRESETn VGND VGND VPWR VPWR _25430_/Q sky130_fd_sc_hd__dfrtp_4
X_22642_ _21058_/A _22641_/X _22303_/X _24872_/Q _22565_/X VGND VGND VPWR VPWR _22643_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_241_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15783__A3 _15782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22573_ _21082_/A _22570_/X _21116_/X _22572_/X VGND VGND VPWR VPWR _22573_/Y sky130_fd_sc_hd__a22oi_4
X_25361_ _25358_/CLK _25361_/D HRESETn VGND VGND VPWR VPWR _25361_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15869__A _21069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24312_ _25543_/CLK _17656_/X HRESETn VGND VGND VPWR VPWR _24312_/Q sky130_fd_sc_hd__dfrtp_4
X_21524_ _21524_/A VGND VGND VPWR VPWR _21524_/Y sky130_fd_sc_hd__inv_2
X_25292_ _25292_/CLK _25292_/D HRESETn VGND VGND VPWR VPWR _11672_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22990__A _21129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21455_ _21042_/X VGND VGND VPWR VPWR _21455_/X sky130_fd_sc_hd__buf_2
X_24243_ _24240_/CLK _18251_/X HRESETn VGND VGND VPWR VPWR _22631_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20406_ _20406_/A VGND VGND VPWR VPWR _20406_/X sky130_fd_sc_hd__buf_2
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24174_ _24201_/CLK _18575_/X HRESETn VGND VGND VPWR VPWR _24174_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21386_ _21386_/A _21386_/B VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__and2_4
XANTENNA__24045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20337_ _21683_/B _20336_/X _20007_/X _20336_/X VGND VGND VPWR VPWR _23430_/D sky130_fd_sc_hd__a2bb2o_4
X_23125_ _16308_/A _23165_/B VGND VGND VPWR VPWR _23125_/X sky130_fd_sc_hd__or2_4
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23056_ _23056_/A _23056_/B VGND VGND VPWR VPWR _23065_/C sky130_fd_sc_hd__and2_4
X_20268_ _20267_/Y _20263_/X _15777_/X _20263_/X VGND VGND VPWR VPWR _20268_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22007_ _22006_/X VGND VGND VPWR VPWR _22007_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20199_ _20197_/Y _20193_/X _20108_/X _20198_/X VGND VGND VPWR VPWR _23482_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12809__B2 _22641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_219_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24537_/CLK sky130_fd_sc_hd__clkbuf_1
X_14760_ _14758_/X _14759_/X _14755_/X VGND VGND VPWR VPWR _25068_/D sky130_fd_sc_hd__o21a_4
XANTENNA__20224__A2_N _20219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11972_ _11967_/A _11660_/A VGND VGND VPWR VPWR _11973_/A sky130_fd_sc_hd__or2_4
X_23958_ _25148_/CLK _23958_/D HRESETn VGND VGND VPWR VPWR _23958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13711_ _11705_/Y _13711_/B VGND VGND VPWR VPWR _13711_/Y sky130_fd_sc_hd__nand2_4
X_22909_ _21090_/A VGND VGND VPWR VPWR _23158_/B sky130_fd_sc_hd__buf_2
XFILLER_204_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14691_ _21275_/A _22085_/A VGND VGND VPWR VPWR _14692_/B sky130_fd_sc_hd__and2_4
X_23889_ _23889_/CLK _19040_/X VGND VGND VPWR VPWR _18090_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_244_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16430_ _16430_/A VGND VGND VPWR VPWR _16430_/Y sky130_fd_sc_hd__inv_2
X_13642_ _13643_/A _13610_/X _13636_/X _13641_/X VGND VGND VPWR VPWR _13642_/X sky130_fd_sc_hd__or4_4
XFILLER_232_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14431__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24886__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _24622_/Q VGND VGND VPWR VPWR _16361_/Y sky130_fd_sc_hd__inv_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12618__D _12618_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13573_ _13565_/X _13567_/X _13573_/C _13573_/D VGND VGND VPWR VPWR _13573_/X sky130_fd_sc_hd__or4_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18155__A _18059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18100_ _18165_/A _18100_/B VGND VGND VPWR VPWR _18100_/X sky130_fd_sc_hd__or2_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19370__B1 _19326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24815__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15312_ _15399_/A _15153_/Y _15423_/A _15396_/A VGND VGND VPWR VPWR _15312_/X sky130_fd_sc_hd__or4_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _25433_/Q VGND VGND VPWR VPWR _12642_/B sky130_fd_sc_hd__inv_2
X_19080_ _19079_/Y _19077_/X _19008_/X _19077_/X VGND VGND VPWR VPWR _19080_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _16287_/Y _16291_/X _11752_/X _16291_/X VGND VGND VPWR VPWR _24648_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18031_ _18031_/A VGND VGND VPWR VPWR _18031_/X sky130_fd_sc_hd__buf_2
X_15243_ _15243_/A _15240_/X VGND VGND VPWR VPWR _15243_/X sky130_fd_sc_hd__or2_4
X_12455_ _12458_/A _12449_/X _12455_/C VGND VGND VPWR VPWR _12455_/X sky130_fd_sc_hd__and3_4
XFILLER_126_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15174_ _15081_/X _15294_/A VGND VGND VPWR VPWR _15174_/X sky130_fd_sc_hd__or2_4
X_12386_ _25346_/Q VGND VGND VPWR VPWR _12386_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14125_ _14125_/A _14125_/B _14111_/A VGND VGND VPWR VPWR _14125_/X sky130_fd_sc_hd__or3_4
XFILLER_125_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19982_ _19981_/Y _19979_/X _19646_/X _19979_/X VGND VGND VPWR VPWR _19982_/X sky130_fd_sc_hd__a2bb2o_4
X_14056_ _14008_/X VGND VGND VPWR VPWR _14056_/Y sky130_fd_sc_hd__inv_2
X_18933_ _18933_/A VGND VGND VPWR VPWR _18933_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21723__A1_N _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13007_ _12999_/X _13052_/B VGND VGND VPWR VPWR _13007_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18864_ _16512_/Y _24145_/Q _16512_/Y _24145_/Q VGND VGND VPWR VPWR _18864_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17815_ _16963_/Y _17815_/B _17814_/X VGND VGND VPWR VPWR _17816_/A sky130_fd_sc_hd__or3_4
X_18795_ _18795_/A VGND VGND VPWR VPWR _18795_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15998__B1 _21091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21108__A1_N _21747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17746_ _17710_/X _17713_/X _17744_/Y _21704_/A _17909_/A VGND VGND VPWR VPWR _17746_/X
+ sky130_fd_sc_hd__a32o_4
X_14958_ _14958_/A VGND VGND VPWR VPWR _14958_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13909_ _13963_/A VGND VGND VPWR VPWR _13954_/B sky130_fd_sc_hd__inv_2
XFILLER_236_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17677_ _17518_/Y _17676_/X VGND VGND VPWR VPWR _17684_/B sky130_fd_sc_hd__or2_4
X_14889_ _14889_/A _14832_/A VGND VGND VPWR VPWR _14889_/Y sky130_fd_sc_hd__nand2_4
XFILLER_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16628_ _16627_/Y _16623_/X _16451_/X _16623_/X VGND VGND VPWR VPWR _24522_/D sky130_fd_sc_hd__a2bb2o_4
X_19416_ _19412_/Y _19415_/X _19326_/X _19415_/X VGND VGND VPWR VPWR _19416_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16559_ _16623_/A VGND VGND VPWR VPWR _16584_/A sky130_fd_sc_hd__buf_2
X_19347_ _19346_/X VGND VGND VPWR VPWR _19353_/A sky130_fd_sc_hd__inv_2
XANTENNA__19361__B1 _19226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12812__A2_N _22726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24556__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19278_ _13757_/C _25282_/Q _13754_/X VGND VGND VPWR VPWR _19278_/X sky130_fd_sc_hd__or3_4
XFILLER_175_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18229_ _18126_/A _19186_/A VGND VGND VPWR VPWR _18229_/X sky130_fd_sc_hd__or2_4
XFILLER_248_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21240_ _21240_/A VGND VGND VPWR VPWR _21273_/A sky130_fd_sc_hd__buf_2
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21171_ _16278_/Y _21574_/A _16192_/A _21170_/X VGND VGND VPWR VPWR _21177_/B sky130_fd_sc_hd__a211o_4
XFILLER_171_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20122_ _20122_/A VGND VGND VPWR VPWR _20122_/X sky130_fd_sc_hd__buf_2
XFILLER_132_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20053_ _20053_/A VGND VGND VPWR VPWR _21477_/B sky130_fd_sc_hd__inv_2
X_24930_ _23678_/CLK _24930_/D HRESETn VGND VGND VPWR VPWR _13603_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_86_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24861_ _24476_/CLK _15780_/X HRESETn VGND VGND VPWR VPWR _24861_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15989__B1 _15632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16650__A1 _15833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23812_ _23628_/CLK _19260_/X VGND VGND VPWR VPWR _23812_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17144__A _17050_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24792_ _24792_/CLK _24792_/D HRESETn VGND VGND VPWR VPWR _21537_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _23735_/CLK _23743_/D VGND VGND VPWR VPWR _18150_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_199_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_192_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24625_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _20954_/X VGND VGND VPWR VPWR _24074_/D sky130_fd_sc_hd__inv_2
XPHY_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_49_0_HCLK clkbuf_7_24_0_HCLK/X VGND VGND VPWR VPWR _24378_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_241_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _23794_/CLK _19661_/X VGND VGND VPWR VPWR _13292_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23279__A2 _22444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20885_/Y _20879_/Y _13671_/B VGND VGND VPWR VPWR _20886_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14413__B1 _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25413_ _24476_/CLK _25413_/D HRESETn VGND VGND VPWR VPWR _12550_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22592_/X _22600_/Y _22625_/C _22624_/Y VGND VGND VPWR VPWR HRDATA[11] sky130_fd_sc_hd__or4_4
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25344_ _25368_/CLK _13114_/Y HRESETn VGND VGND VPWR VPWR _12372_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22556_ _22555_/X VGND VGND VPWR VPWR _22556_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21507_ _21815_/A _21505_/X _21507_/C VGND VGND VPWR VPWR _21507_/X sky130_fd_sc_hd__and3_4
X_25275_ _25103_/CLK _13832_/X HRESETn VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15913__B1 _15636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22487_ _22487_/A _22486_/X VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__and2_4
X_12240_ _21451_/A VGND VGND VPWR VPWR _12240_/Y sky130_fd_sc_hd__inv_2
X_24226_ _24230_/CLK _24226_/D HRESETn VGND VGND VPWR VPWR _23360_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22870__D _22869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21438_ _21431_/X _21432_/X _21434_/X _24861_/Q _22558_/A VGND VGND VPWR VPWR _21439_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12171_ _14342_/B VGND VGND VPWR VPWR _12172_/B sky130_fd_sc_hd__inv_2
XFILLER_135_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21369_ _21369_/A _21369_/B VGND VGND VPWR VPWR _21369_/Y sky130_fd_sc_hd__nand2_4
X_24157_ _24160_/CLK _18732_/Y HRESETn VGND VGND VPWR VPWR _24157_/Q sky130_fd_sc_hd__dfrtp_4
X_23108_ _16115_/Y _22569_/X _22861_/X _11775_/Y _22864_/X VGND VGND VPWR VPWR _23108_/X
+ sky130_fd_sc_hd__o32a_4
X_24088_ _23980_/CLK _20522_/X HRESETn VGND VGND VPWR VPWR _24088_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15930_ _15694_/X _15928_/Y _15686_/X _15928_/Y VGND VGND VPWR VPWR _15930_/X sky130_fd_sc_hd__a2bb2o_4
X_23039_ _16733_/A _23036_/X _23038_/X VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__and3_4
XANTENNA__25085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17969__A1 _18069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17969__B2 _15694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15861_ _21592_/A VGND VGND VPWR VPWR _21589_/B sky130_fd_sc_hd__buf_2
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17600_ _17895_/B VGND VGND VPWR VPWR _17600_/X sky130_fd_sc_hd__buf_2
XFILLER_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14812_ _14826_/C _14811_/X _14812_/C VGND VGND VPWR VPWR _14812_/X sky130_fd_sc_hd__or3_4
XFILLER_18_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18580_ _18476_/B _18570_/X VGND VGND VPWR VPWR _18581_/C sky130_fd_sc_hd__nand2_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15792_ _15792_/A VGND VGND VPWR VPWR _15792_/X sky130_fd_sc_hd__buf_2
XANTENNA__22895__A _23008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14901__A2_N _14899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17531_ _17531_/A VGND VGND VPWR VPWR _17531_/Y sky130_fd_sc_hd__inv_2
X_14743_ _25073_/Q VGND VGND VPWR VPWR _22060_/A sky130_fd_sc_hd__inv_2
XANTENNA__17989__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11955_ _19643_/A VGND VGND VPWR VPWR _11955_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17462_ _13182_/A _17461_/X VGND VGND VPWR VPWR _17466_/A sky130_fd_sc_hd__and2_4
X_14674_ _14674_/A VGND VGND VPWR VPWR _14674_/X sky130_fd_sc_hd__buf_2
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11886_ _11886_/A _11885_/X VGND VGND VPWR VPWR _11887_/B sky130_fd_sc_hd__and2_4
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16413_ _15156_/Y _16409_/X _16412_/X _16409_/X VGND VGND VPWR VPWR _24605_/D sky130_fd_sc_hd__a2bb2o_4
X_19201_ _19200_/Y _19196_/X _19131_/X _19196_/X VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13625_ _18102_/A VGND VGND VPWR VPWR _13625_/X sky130_fd_sc_hd__buf_2
XANTENNA__21304__A _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17393_ _17251_/A _17393_/B VGND VGND VPWR VPWR _17393_/X sky130_fd_sc_hd__or2_4
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19132_ _19130_/Y _19126_/X _19131_/X _19126_/X VGND VGND VPWR VPWR _19132_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11830__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16344_ _16343_/Y _16339_/X _16248_/X _16339_/X VGND VGND VPWR VPWR _24629_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13556_ _13555_/Y _14567_/A _13555_/Y _14567_/A VGND VGND VPWR VPWR _13556_/X sky130_fd_sc_hd__a2bb2o_4
X_12507_ _12513_/A _12478_/B VGND VGND VPWR VPWR _12514_/B sky130_fd_sc_hd__or2_4
X_19063_ _23881_/Q VGND VGND VPWR VPWR _19063_/Y sky130_fd_sc_hd__inv_2
X_16275_ _21340_/A VGND VGND VPWR VPWR _16275_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15021__B _15021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13487_ _13483_/Y _13486_/X _11842_/X _13486_/X VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_139_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18014_ _18200_/A _23899_/Q VGND VGND VPWR VPWR _18015_/C sky130_fd_sc_hd__or2_4
X_15226_ _15075_/D _15220_/X _15208_/X _15223_/B VGND VGND VPWR VPWR _15227_/A sky130_fd_sc_hd__a211o_4
X_12438_ _12514_/A VGND VGND VPWR VPWR _12458_/A sky130_fd_sc_hd__buf_2
XANTENNA__21453__A1 _21307_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15157_ _15096_/Y _24611_/Q _25001_/Q _15156_/Y VGND VGND VPWR VPWR _15161_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21453__B2 _22531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20116__A2_N _20109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12369_ _12362_/X _12369_/B _12369_/C _12369_/D VGND VGND VPWR VPWR _12390_/B sky130_fd_sc_hd__or4_4
XFILLER_154_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14108_ _25219_/Q _14108_/B _14108_/C VGND VGND VPWR VPWR _14109_/B sky130_fd_sc_hd__or3_4
X_15088_ _24987_/Q _15086_/Y _15340_/A _15099_/A VGND VGND VPWR VPWR _15091_/C sky130_fd_sc_hd__a2bb2o_4
X_19965_ _19965_/A _19480_/X _19505_/X VGND VGND VPWR VPWR _19965_/X sky130_fd_sc_hd__or3_4
XANTENNA__22789__B _22789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15972__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14039_ _14037_/Y _14039_/B _14010_/X _14022_/A VGND VGND VPWR VPWR _14040_/A sky130_fd_sc_hd__or4_4
X_18916_ _18916_/A VGND VGND VPWR VPWR _18916_/Y sky130_fd_sc_hd__inv_2
X_19896_ _19894_/Y _19895_/X _19643_/X _19895_/X VGND VGND VPWR VPWR _23591_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14891__B1 _14890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24005__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ _24579_/Q _18703_/A _16546_/Y _24132_/Q VGND VGND VPWR VPWR _18850_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18778_ _18777_/X VGND VGND VPWR VPWR _24145_/D sky130_fd_sc_hd__inv_2
XFILLER_243_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18909__B1 _18908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_202_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _24194_/CLK sky130_fd_sc_hd__clkbuf_1
X_17729_ _24219_/Q VGND VGND VPWR VPWR _17729_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13642__D _13641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24737__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_8_0_HCLK clkbuf_8_9_0_HCLK/A VGND VGND VPWR VPWR _23563_/CLK sky130_fd_sc_hd__clkbuf_1
X_20740_ _13139_/X VGND VGND VPWR VPWR _20740_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16396__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20671_ _20670_/X VGND VGND VPWR VPWR _23997_/D sky130_fd_sc_hd__inv_2
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19334__B1 _19220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _21288_/X _22406_/Y _21525_/Y _22409_/X VGND VGND VPWR VPWR _22410_/X sky130_fd_sc_hd__a2bb2o_4
X_23390_ _23913_/CLK _23390_/D VGND VGND VPWR VPWR _13353_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22341_ _22334_/Y _22336_/Y _22337_/X _22340_/Y _21565_/Y VGND VGND VPWR VPWR _22341_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21868__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22272_ _21472_/A _22272_/B _22272_/C VGND VGND VPWR VPWR _22272_/X sky130_fd_sc_hd__and3_4
X_25060_ _23385_/CLK _25060_/D HRESETn VGND VGND VPWR VPWR _14806_/A sky130_fd_sc_hd__dfrtp_4
X_21223_ _13789_/X _21221_/X _22527_/A _21222_/X VGND VGND VPWR VPWR _21224_/A sky130_fd_sc_hd__a211o_4
X_24011_ _25106_/CLK _20468_/X HRESETn VGND VGND VPWR VPWR _24011_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21154_ _12132_/Y _21031_/X _21583_/B _21153_/Y VGND VGND VPWR VPWR _21154_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21884__A _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20105_ _20105_/A VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__buf_2
X_21085_ _21085_/A VGND VGND VPWR VPWR _21085_/X sky130_fd_sc_hd__buf_2
XFILLER_101_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20036_ _23540_/Q VGND VGND VPWR VPWR _22347_/B sky130_fd_sc_hd__inv_2
X_24913_ _24913_/CLK _15610_/X HRESETn VGND VGND VPWR VPWR _15608_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24844_ _25425_/CLK _15822_/X HRESETn VGND VGND VPWR VPWR _24844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15001__A2_N _24452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24775_ _24777_/CLK _24775_/D HRESETn VGND VGND VPWR VPWR _24775_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ _20413_/Y _21972_/B VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__or2_4
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A _13786_/A _11740_/C _11740_/D VGND VGND VPWR VPWR _15661_/C sky130_fd_sc_hd__or4_4
X_23726_ _23717_/CLK _19499_/X VGND VGND VPWR VPWR _23726_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _16671_/Y _20854_/A _20863_/X _20937_/X VGND VGND VPWR VPWR _20939_/A sky130_fd_sc_hd__o22a_4
XFILLER_230_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11672_/A _11670_/Y _13693_/A _24235_/Q VGND VGND VPWR VPWR _11675_/C sky130_fd_sc_hd__a2bb2o_4
X_23657_ _23642_/CLK _19707_/X VGND VGND VPWR VPWR _13326_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20824__A1_N _20698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _24055_/Q VGND VGND VPWR VPWR _20870_/C sky130_fd_sc_hd__inv_2
XFILLER_202_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13410_/A _23870_/Q VGND VGND VPWR VPWR _13412_/B sky130_fd_sc_hd__or2_4
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22608_ _22608_/A _21450_/X VGND VGND VPWR VPWR _22608_/X sky130_fd_sc_hd__or2_4
XANTENNA__16139__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14390_ _14116_/A _14390_/B VGND VGND VPWR VPWR _14392_/A sky130_fd_sc_hd__nor2_4
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23588_ _23684_/CLK _23588_/D VGND VGND VPWR VPWR _23588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13332_/X _13335_/X _13340_/X VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__or3_4
X_25327_ _25181_/CLK _25327_/D HRESETn VGND VGND VPWR VPWR _13490_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22539_ _23313_/B VGND VGND VPWR VPWR _22589_/B sky130_fd_sc_hd__buf_2
XFILLER_127_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16060_ _24730_/Q VGND VGND VPWR VPWR _16060_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13272_ _13411_/A _13272_/B VGND VGND VPWR VPWR _13273_/C sky130_fd_sc_hd__or2_4
X_25258_ _25204_/CLK _13868_/X HRESETn VGND VGND VPWR VPWR _25258_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15901__A3 _16248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15011_ _15011_/A _15011_/B _15011_/C _15010_/X VGND VGND VPWR VPWR _15011_/X sky130_fd_sc_hd__or4_4
X_12223_ _22910_/A VGND VGND VPWR VPWR _12223_/Y sky130_fd_sc_hd__inv_2
X_24209_ _24111_/CLK _18353_/X HRESETn VGND VGND VPWR VPWR _13211_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22632__B1 _21968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25189_ _23385_/CLK _25189_/D HRESETn VGND VGND VPWR VPWR _25189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12154_ _12144_/X _12145_/X _12149_/X _12153_/X VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__or4_4
X_19750_ _19750_/A VGND VGND VPWR VPWR _19750_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19264__A _19258_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12085_ _12085_/A VGND VGND VPWR VPWR _12085_/Y sky130_fd_sc_hd__inv_2
X_16962_ _16962_/A _16961_/X VGND VGND VPWR VPWR _16962_/X sky130_fd_sc_hd__or2_4
XFILLER_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18701_ _18701_/A _18733_/A _18701_/C _18733_/B VGND VGND VPWR VPWR _18701_/X sky130_fd_sc_hd__or4_4
X_15913_ _12805_/Y _15912_/X _15636_/X _15912_/X VGND VGND VPWR VPWR _24795_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16893_ _19810_/A VGND VGND VPWR VPWR _16893_/Y sky130_fd_sc_hd__inv_2
X_19681_ _19681_/A VGND VGND VPWR VPWR _19681_/Y sky130_fd_sc_hd__inv_2
X_15844_ _15844_/A VGND VGND VPWR VPWR _15844_/X sky130_fd_sc_hd__buf_2
X_18632_ _18632_/A _18627_/X _18629_/X _18631_/X VGND VGND VPWR VPWR _18632_/X sky130_fd_sc_hd__or4_4
XFILLER_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14201__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15775_ _11855_/A VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__buf_2
X_18563_ _18484_/B _18558_/B _18560_/B _18494_/X VGND VGND VPWR VPWR _18564_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22699__B1 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12987_ _21035_/A _12640_/B VGND VGND VPWR VPWR _12988_/C sky130_fd_sc_hd__or2_4
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24830__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14726_ _13744_/A _13768_/A _25285_/Q _13768_/Y VGND VGND VPWR VPWR _14726_/X sky130_fd_sc_hd__o22a_4
X_17514_ _11873_/Y _24296_/Q _11873_/Y _24296_/Q VGND VGND VPWR VPWR _17515_/D sky130_fd_sc_hd__a2bb2o_4
X_11938_ _19629_/A VGND VGND VPWR VPWR _11938_/Y sky130_fd_sc_hd__inv_2
X_18494_ _18828_/B VGND VGND VPWR VPWR _18494_/X sky130_fd_sc_hd__buf_2
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17445_ _17445_/A VGND VGND VPWR VPWR _17445_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21034__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14657_ _18130_/A VGND VGND VPWR VPWR _17945_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_32_0_HCLK clkbuf_8_33_0_HCLK/A VGND VGND VPWR VPWR _23577_/CLK sky130_fd_sc_hd__clkbuf_1
X_11869_ _11869_/A VGND VGND VPWR VPWR _11869_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_95_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _25433_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ _14679_/B VGND VGND VPWR VPWR _14668_/A sky130_fd_sc_hd__buf_2
X_17376_ _17198_/X _17375_/X _17280_/X VGND VGND VPWR VPWR _17376_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14588_ _14593_/A _14582_/Y VGND VGND VPWR VPWR _14588_/X sky130_fd_sc_hd__and2_4
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16327_ _24635_/Q VGND VGND VPWR VPWR _16327_/Y sky130_fd_sc_hd__inv_2
X_19115_ _21400_/B _19112_/X _16897_/X _19112_/X VGND VGND VPWR VPWR _23862_/D sky130_fd_sc_hd__a2bb2o_4
X_13539_ _13526_/Y _13538_/Y SCLK_S2 _13537_/X VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__o22a_4
XFILLER_173_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17878__B1 _16964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15967__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19046_ _18189_/B VGND VGND VPWR VPWR _19046_/Y sky130_fd_sc_hd__inv_2
X_16258_ _16256_/Y _16251_/X _16153_/X _16257_/X VGND VGND VPWR VPWR _24661_/D sky130_fd_sc_hd__a2bb2o_4
X_15209_ _15203_/A _15202_/X _15208_/X _15204_/Y VGND VGND VPWR VPWR _15210_/A sky130_fd_sc_hd__a211o_4
XFILLER_127_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16189_ _23341_/A VGND VGND VPWR VPWR _16189_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19174__A _19181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19948_ _19948_/A VGND VGND VPWR VPWR _22264_/B sky130_fd_sc_hd__inv_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22312__B _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19879_ _19878_/Y _19874_/X _19856_/X _19861_/Y VGND VGND VPWR VPWR _23597_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21910_ _22094_/A _21910_/B VGND VGND VPWR VPWR _21911_/C sky130_fd_sc_hd__or2_4
XANTENNA__11735__A _21135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22890_ _16684_/Y _22890_/B VGND VGND VPWR VPWR _22890_/X sky130_fd_sc_hd__and2_4
XANTENNA__18070__A3 _18069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15959__A3 HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18651__A1_N _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21841_ _21841_/A _21762_/X _21841_/C _21840_/X VGND VGND VPWR VPWR HRDATA[3] sky130_fd_sc_hd__or4_4
XFILLER_209_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21870__C _21752_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19555__B1 _19418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24571__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17422__A _17422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24560_ _24528_/CLK _16528_/X HRESETn VGND VGND VPWR VPWR _24560_/Q sky130_fd_sc_hd__dfrtp_4
X_21772_ _21646_/A _21770_/X _21771_/X VGND VGND VPWR VPWR _21772_/X sky130_fd_sc_hd__and3_4
XANTENNA__16369__B1 _16368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21362__B1 SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _24295_/CLK _23511_/D VGND VGND VPWR VPWR _23511_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22928__A1_N _17263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20723_ _20722_/X VGND VGND VPWR VPWR _24021_/D sky130_fd_sc_hd__inv_2
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24491_ _24666_/CLK _16712_/X HRESETn VGND VGND VPWR VPWR _24491_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18666__A1_N _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23555_/CLK _23442_/D VGND VGND VPWR VPWR _20305_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21879__A _21879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20654_ _14250_/Y _20646_/X _20637_/X _20653_/X VGND VGND VPWR VPWR _20654_/X sky130_fd_sc_hd__a211o_4
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_3_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20585_ _20588_/B _20584_/Y _20597_/C VGND VGND VPWR VPWR _20585_/X sky130_fd_sc_hd__and3_4
X_23373_ _23360_/X VGND VGND VPWR VPWR IRQ[17] sky130_fd_sc_hd__buf_2
X_25112_ _23970_/CLK _25112_/D HRESETn VGND VGND VPWR VPWR _25112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22324_ _23937_/Q VGND VGND VPWR VPWR _22324_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16541__B1 _16364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25043_ _25043_/CLK _25043_/D HRESETn VGND VGND VPWR VPWR _25043_/Q sky130_fd_sc_hd__dfrtp_4
X_22255_ _22260_/A _22255_/B VGND VGND VPWR VPWR _22257_/B sky130_fd_sc_hd__or2_4
XFILLER_164_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21206_ _21204_/A VGND VGND VPWR VPWR _21209_/A sky130_fd_sc_hd__buf_2
X_22186_ _13512_/Y _12107_/A _12040_/Y _12080_/A VGND VGND VPWR VPWR _22186_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22503__A _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21137_ _25107_/Q _21351_/A VGND VGND VPWR VPWR _21143_/A sky130_fd_sc_hd__nand2_4
XFILLER_87_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21068_ _22533_/A VGND VGND VPWR VPWR _21068_/X sky130_fd_sc_hd__buf_2
XFILLER_219_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23037__C _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24659__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12988_/A VGND VGND VPWR VPWR _12927_/A sky130_fd_sc_hd__buf_2
X_20019_ _23547_/Q VGND VGND VPWR VPWR _20019_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13890_ _13880_/X _13889_/X _25191_/Q _13876_/A VGND VGND VPWR VPWR _13890_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12841_ _25401_/Q _12829_/Y _12828_/X _24794_/Q VGND VGND VPWR VPWR _12844_/C sky130_fd_sc_hd__a2bb2o_4
X_24827_ _24849_/CLK _15847_/X HRESETn VGND VGND VPWR VPWR _24827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15560_ _14386_/A _21122_/A VGND VGND VPWR VPWR _15560_/X sky130_fd_sc_hd__or2_4
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12772_ _12772_/A _12766_/X _12772_/C _12771_/X VGND VGND VPWR VPWR _12772_/X sky130_fd_sc_hd__or4_4
X_24758_ _24767_/CLK _15991_/X HRESETn VGND VGND VPWR VPWR _22159_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16959__A2_N _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _23969_/Q VGND VGND VPWR VPWR _14524_/A sky130_fd_sc_hd__buf_2
XFILLER_214_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _24079_/Q VGND VGND VPWR VPWR _11724_/A sky130_fd_sc_hd__inv_2
X_23709_ _23717_/CLK _23709_/D VGND VGND VPWR VPWR _23709_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _24955_/Q _15447_/X _15444_/X VGND VGND VPWR VPWR _24955_/D sky130_fd_sc_hd__a21bo_4
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24689_/CLK _24689_/D HRESETn VGND VGND VPWR VPWR _21709_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _16304_/Y _17245_/A _16322_/A _17229_/Y VGND VGND VPWR VPWR _17233_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A VGND VGND VPWR VPWR _14443_/A sky130_fd_sc_hd__buf_2
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21789__A _22387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16780__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22448__A3 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19849__B2 _19844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _17051_/Y _17138_/B _17159_/B _17076_/X VGND VGND VPWR VPWR _17162_/A sky130_fd_sc_hd__a211o_4
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _25163_/Q _14360_/X _25162_/Q _14365_/X VGND VGND VPWR VPWR _14373_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19259__A _19258_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _16110_/Y _16111_/X _11770_/X _16111_/X VGND VGND VPWR VPWR _16112_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13456_/A _13315_/X _13324_/C VGND VGND VPWR VPWR _13324_/X sky130_fd_sc_hd__and3_4
X_17092_ _17095_/A _17088_/X _17091_/Y VGND VGND VPWR VPWR _17092_/X sky130_fd_sc_hd__and3_4
XFILLER_171_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16043_ _16004_/X VGND VGND VPWR VPWR _16044_/A sky130_fd_sc_hd__buf_2
X_13255_ _13155_/X VGND VGND VPWR VPWR _13428_/A sky130_fd_sc_hd__buf_2
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12206_ _12205_/Y _21091_/A _12205_/Y _21091_/A VGND VGND VPWR VPWR _12206_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13186_ _13306_/A VGND VGND VPWR VPWR _13186_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19802_ _19802_/A VGND VGND VPWR VPWR _21766_/B sky130_fd_sc_hd__inv_2
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12137_ _24117_/Q _12150_/A VGND VGND VPWR VPWR _12138_/A sky130_fd_sc_hd__and2_4
XFILLER_150_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17994_ _17985_/A VGND VGND VPWR VPWR _18178_/A sky130_fd_sc_hd__buf_2
XANTENNA__13527__A1_N _13526_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19733_ _19719_/Y VGND VGND VPWR VPWR _19733_/X sky130_fd_sc_hd__buf_2
XANTENNA__23030__B1 _16952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12068_ _17448_/C VGND VGND VPWR VPWR _12068_/X sky130_fd_sc_hd__buf_2
X_16945_ _16138_/Y _17764_/A _16138_/Y _17764_/A VGND VGND VPWR VPWR _16945_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19785__B1 _19761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12321__B2 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19664_ _13365_/B VGND VGND VPWR VPWR _19664_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16876_ _16870_/X VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__buf_2
XFILLER_231_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18615_ _18614_/Y VGND VGND VPWR VPWR _18794_/C sky130_fd_sc_hd__buf_2
X_15827_ _15825_/X _15804_/X _15748_/X _24841_/Q _15826_/X VGND VGND VPWR VPWR _15827_/X
+ sky130_fd_sc_hd__a32o_4
X_19595_ _19595_/A _21161_/A VGND VGND VPWR VPWR _21380_/A sky130_fd_sc_hd__or2_4
XFILLER_231_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22136__A2 _22119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ _15758_/A VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__buf_2
X_18546_ _18550_/A _18540_/X _18546_/C VGND VGND VPWR VPWR _18546_/X sky130_fd_sc_hd__and3_4
XFILLER_178_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14709_ _21262_/A VGND VGND VPWR VPWR _14709_/X sky130_fd_sc_hd__buf_2
XANTENNA__11832__B1 _11831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15689_ _24893_/Q VGND VGND VPWR VPWR _15696_/A sky130_fd_sc_hd__inv_2
X_18477_ _24166_/Q VGND VGND VPWR VPWR _18595_/A sky130_fd_sc_hd__inv_2
XFILLER_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17428_ _20680_/A _17426_/X _17427_/X _17426_/X VGND VGND VPWR VPWR _17428_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21699__A _22274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16771__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12388__B2 _24828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _17364_/A _17364_/B _17359_/C _17364_/C VGND VGND VPWR VPWR _17360_/A sky130_fd_sc_hd__or4_4
XANTENNA__25188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20370_ _20364_/Y VGND VGND VPWR VPWR _20370_/X sky130_fd_sc_hd__buf_2
XFILLER_174_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16523__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19029_ _19028_/X VGND VGND VPWR VPWR _19037_/A sky130_fd_sc_hd__inv_2
X_22040_ _22029_/A _22038_/X _22040_/C VGND VGND VPWR VPWR _22040_/X sky130_fd_sc_hd__and3_4
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23991_ _23991_/CLK _23991_/D HRESETn VGND VGND VPWR VPWR _17400_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19776__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24752__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22942_ _24571_/Q _22897_/X _22816_/X VGND VGND VPWR VPWR _22942_/X sky130_fd_sc_hd__o21a_4
XFILLER_217_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24124__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22873_ _22777_/X _22871_/X _22872_/X _24843_/Q _22779_/X VGND VGND VPWR VPWR _22873_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24612_ _24602_/CLK _24612_/D HRESETn VGND VGND VPWR VPWR _15099_/A sky130_fd_sc_hd__dfrtp_4
X_21824_ _21820_/X _21823_/X _21499_/X VGND VGND VPWR VPWR _21832_/B sky130_fd_sc_hd__o21a_4
XFILLER_231_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24543_ _24542_/CLK _24543_/D HRESETn VGND VGND VPWR VPWR _16574_/A sky130_fd_sc_hd__dfrtp_4
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21886__A1 _16166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11823__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21755_ _21755_/A _21755_/B VGND VGND VPWR VPWR _21762_/C sky130_fd_sc_hd__nor2_4
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21886__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _15643_/Y _20695_/X _20704_/X _20705_/X VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__o22a_4
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _24473_/CLK _16755_/X HRESETn VGND VGND VPWR VPWR _16754_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21686_ _21685_/X VGND VGND VPWR VPWR _22029_/A sky130_fd_sc_hd__buf_2
XFILLER_212_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23425_ _23493_/CLK _23425_/D VGND VGND VPWR VPWR _21996_/C sky130_fd_sc_hd__dfxtp_4
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20637_ _20637_/A VGND VGND VPWR VPWR _20637_/X sky130_fd_sc_hd__buf_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23356_ _25276_/Q _23356_/B VGND VGND VPWR VPWR _23356_/X sky130_fd_sc_hd__and2_4
XANTENNA__16514__B1 _16241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20568_ _14450_/Y _20551_/X _20565_/X _20567_/X VGND VGND VPWR VPWR _20569_/A sky130_fd_sc_hd__a211o_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22307_ _13667_/A VGND VGND VPWR VPWR _22307_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23287_ _24783_/Q _22669_/B VGND VGND VPWR VPWR _23287_/X sky130_fd_sc_hd__or2_4
XFILLER_164_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20499_ _23978_/Q _20487_/B _20499_/C VGND VGND VPWR VPWR _20499_/X sky130_fd_sc_hd__and3_4
XFILLER_166_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13040_ _13049_/A VGND VGND VPWR VPWR _13040_/X sky130_fd_sc_hd__buf_2
X_25026_ _25023_/CLK _15252_/X HRESETn VGND VGND VPWR VPWR _15250_/A sky130_fd_sc_hd__dfrtp_4
X_22238_ _21981_/B _19597_/X VGND VGND VPWR VPWR _22238_/X sky130_fd_sc_hd__and2_4
XFILLER_180_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22169_ _15037_/A _21312_/B _21335_/X VGND VGND VPWR VPWR _22169_/X sky130_fd_sc_hd__o21a_4
XFILLER_121_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14991_ _15276_/A _24425_/Q _14990_/X _24422_/Q VGND VGND VPWR VPWR _14991_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13942_ _13942_/A VGND VGND VPWR VPWR _13942_/X sky130_fd_sc_hd__buf_2
X_16730_ _16728_/Y _16654_/X _16729_/X _16654_/X VGND VGND VPWR VPWR _24484_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12597__A2_N _12595_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16661_ _23244_/A _16655_/X _16393_/X _16660_/X VGND VGND VPWR VPWR _24512_/D sky130_fd_sc_hd__a2bb2o_4
X_13873_ _13871_/A _13870_/X _13871_/Y _13872_/X VGND VGND VPWR VPWR _13873_/X sky130_fd_sc_hd__o22a_4
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15253__B1 _15208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15612_ _15611_/Y _15609_/X _11813_/X _15609_/X VGND VGND VPWR VPWR _24912_/D sky130_fd_sc_hd__a2bb2o_4
X_18400_ _24169_/Q VGND VGND VPWR VPWR _18400_/Y sky130_fd_sc_hd__inv_2
X_12824_ _12824_/A _12824_/B _12824_/C _12823_/X VGND VGND VPWR VPWR _12845_/B sky130_fd_sc_hd__or4_4
X_16592_ _16618_/A VGND VGND VPWR VPWR _16592_/X sky130_fd_sc_hd__buf_2
X_19380_ _19379_/Y _19374_/X _19246_/X _19374_/X VGND VGND VPWR VPWR _23768_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15543_ _16462_/C _15538_/X HADDR[5] _15538_/X VGND VGND VPWR VPWR _15543_/X sky130_fd_sc_hd__a2bb2o_4
X_18331_ _24213_/Q VGND VGND VPWR VPWR _18959_/A sky130_fd_sc_hd__buf_2
XFILLER_43_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12755_ _22302_/A VGND VGND VPWR VPWR _12755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17997__A _18102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12520__A2_N _24871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _24244_/Q VGND VGND VPWR VPWR _11706_/Y sky130_fd_sc_hd__inv_2
X_18262_ _20408_/A VGND VGND VPWR VPWR _18262_/X sky130_fd_sc_hd__buf_2
XFILLER_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _24962_/Q VGND VGND VPWR VPWR _15474_/Y sky130_fd_sc_hd__inv_2
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12618_/A _12691_/B _12662_/X VGND VGND VPWR VPWR _12686_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16753__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14425_/A VGND VGND VPWR VPWR _14425_/Y sky130_fd_sc_hd__inv_2
X_17213_ _24634_/Q _17330_/A _16361_/Y _24351_/Q VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18193_ _18129_/A _19022_/A VGND VGND VPWR VPWR _18194_/C sky130_fd_sc_hd__or2_4
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_106_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24629_/CLK sky130_fd_sc_hd__clkbuf_1
X_17144_ _17050_/D _17143_/X VGND VGND VPWR VPWR _17144_/X sky130_fd_sc_hd__or2_4
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14349_/A _14359_/B _14355_/Y VGND VGND VPWR VPWR _25169_/D sky130_fd_sc_hd__o21a_4
XFILLER_11_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16505__B1 _16419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_169_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23880_/CLK sky130_fd_sc_hd__clkbuf_1
X_13307_ _13417_/A _13307_/B VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__or2_4
X_17075_ _17035_/Y _17057_/X _17075_/C _17074_/X VGND VGND VPWR VPWR _17075_/X sky130_fd_sc_hd__or4_4
X_14287_ _14286_/Y VGND VGND VPWR VPWR _15465_/A sky130_fd_sc_hd__buf_2
XFILLER_170_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16026_ _24744_/Q VGND VGND VPWR VPWR _16026_/Y sky130_fd_sc_hd__inv_2
X_13238_ _13322_/A _13238_/B _13237_/X VGND VGND VPWR VPWR _13239_/C sky130_fd_sc_hd__and3_4
XFILLER_170_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22143__A _21300_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13169_ _13197_/A _13169_/B _13168_/X VGND VGND VPWR VPWR _13169_/X sky130_fd_sc_hd__and3_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17977_ _17977_/A _23771_/Q VGND VGND VPWR VPWR _17977_/X sky130_fd_sc_hd__or2_4
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19716_ _19715_/Y _19711_/X _19620_/X _19698_/Y VGND VGND VPWR VPWR _19716_/X sky130_fd_sc_hd__a2bb2o_4
X_16928_ _22502_/A _17871_/A _16152_/Y _17861_/A VGND VGND VPWR VPWR _16928_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19647_ _21506_/B _19642_/X _19646_/X _19642_/X VGND VGND VPWR VPWR _19647_/X sky130_fd_sc_hd__a2bb2o_4
X_16859_ _24422_/Q VGND VGND VPWR VPWR _16859_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22109__A2 _21069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19578_ _22247_/B _19575_/X _11943_/X _19575_/X VGND VGND VPWR VPWR _23699_/D sky130_fd_sc_hd__a2bb2o_4
X_18529_ _18515_/A _18515_/B VGND VGND VPWR VPWR _18538_/B sky130_fd_sc_hd__or2_4
XANTENNA__25369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _21714_/A _21540_/B VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__and2_4
XANTENNA__16744__B1 _16389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21222__A _24328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22817__B1 _22816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21471_ _21209_/A VGND VGND VPWR VPWR _21472_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_65_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23210_ _17294_/A _22493_/X _12888_/A _22453_/X VGND VGND VPWR VPWR _23210_/X sky130_fd_sc_hd__a2bb2o_4
X_20422_ _20422_/A VGND VGND VPWR VPWR _20422_/Y sky130_fd_sc_hd__inv_2
X_24190_ _24194_/CLK _18511_/X HRESETn VGND VGND VPWR VPWR _24190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23141_ _23137_/X _23138_/X _23139_/X _23140_/X VGND VGND VPWR VPWR _23142_/B sky130_fd_sc_hd__o22a_4
XFILLER_146_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20353_ _20350_/Y _20352_/X _20243_/X _20352_/X VGND VGND VPWR VPWR _23424_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20284_ _20278_/Y VGND VGND VPWR VPWR _20284_/X sky130_fd_sc_hd__buf_2
X_23072_ _23072_/A _23072_/B VGND VGND VPWR VPWR _23072_/Y sky130_fd_sc_hd__nor2_4
XFILLER_1_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23242__B1 _25401_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22023_ _22027_/A VGND VGND VPWR VPWR _22032_/A sky130_fd_sc_hd__buf_2
XFILLER_121_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17147__A _17050_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_25_0_HCLK_A clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23974_ _23976_/CLK _23974_/D HRESETn VGND VGND VPWR VPWR _23974_/Q sky130_fd_sc_hd__dfrtp_4
X_22925_ _12222_/Y _22507_/X _24282_/Q _22924_/X VGND VGND VPWR VPWR _22930_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22856_ _16733_/A _22856_/B _22855_/X VGND VGND VPWR VPWR _22856_/X sky130_fd_sc_hd__and3_4
X_21807_ _21673_/A _21807_/B VGND VGND VPWR VPWR _21807_/X sky130_fd_sc_hd__or2_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18925__A2_N _18922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22787_ _22437_/X VGND VGND VPWR VPWR _22787_/X sky130_fd_sc_hd__buf_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12540_ _12531_/X _12534_/X _12537_/X _12540_/D VGND VGND VPWR VPWR _12540_/X sky130_fd_sc_hd__or4_4
X_24526_ _24528_/CLK _24526_/D HRESETn VGND VGND VPWR VPWR _16617_/A sky130_fd_sc_hd__dfrtp_4
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21738_ _21738_/A VGND VGND VPWR VPWR _21739_/D sky130_fd_sc_hd__inv_2
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16735__B1 _16729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21132__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12471_ _12250_/A _12470_/Y VGND VGND VPWR VPWR _12473_/B sky130_fd_sc_hd__or2_4
X_24457_ _24425_/CLK _16788_/X HRESETn VGND VGND VPWR VPWR _15037_/A sky130_fd_sc_hd__dfrtp_4
X_21669_ _21673_/A _20050_/Y VGND VGND VPWR VPWR _21669_/X sky130_fd_sc_hd__or2_4
XFILLER_200_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14210_ _14210_/A VGND VGND VPWR VPWR _14210_/X sky130_fd_sc_hd__buf_2
X_23408_ _23408_/CLK _23408_/D VGND VGND VPWR VPWR _23408_/Q sky130_fd_sc_hd__dfxtp_4
X_15190_ _15068_/X _15190_/B _15190_/C VGND VGND VPWR VPWR _15190_/X sky130_fd_sc_hd__and3_4
XFILLER_172_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24388_ _24386_/CLK _17148_/X HRESETn VGND VGND VPWR VPWR _16974_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14141_ _14141_/A VGND VGND VPWR VPWR _23967_/D sky130_fd_sc_hd__buf_2
X_23339_ _13147_/A _21296_/X _13677_/A _21320_/X VGND VGND VPWR VPWR _23339_/Y sky130_fd_sc_hd__a22oi_4
X_14072_ _20470_/B VGND VGND VPWR VPWR _14073_/A sky130_fd_sc_hd__buf_2
X_13023_ _13023_/A _13022_/Y VGND VGND VPWR VPWR _13025_/B sky130_fd_sc_hd__or2_4
X_17900_ _17900_/A VGND VGND VPWR VPWR _17900_/Y sky130_fd_sc_hd__inv_2
X_25009_ _25002_/CLK _15336_/Y HRESETn VGND VGND VPWR VPWR _25009_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24674__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18880_ _20570_/A _20567_/A VGND VGND VPWR VPWR _20571_/A sky130_fd_sc_hd__or2_4
XANTENNA__18255__A3 _16609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21795__B1 _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24603__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17831_ _17768_/D _17820_/B VGND VGND VPWR VPWR _17832_/B sky130_fd_sc_hd__or2_4
XFILLER_79_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18660__B1 _16606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17762_ _17762_/A VGND VGND VPWR VPWR _17762_/Y sky130_fd_sc_hd__inv_2
X_14974_ _14973_/Y _14980_/A _25023_/Q _14909_/Y VGND VGND VPWR VPWR _14983_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_248_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19501_ _19900_/A VGND VGND VPWR VPWR _19501_/X sky130_fd_sc_hd__buf_2
X_16713_ _16713_/A VGND VGND VPWR VPWR _16713_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21307__A _24485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13925_ _13924_/X VGND VGND VPWR VPWR _14260_/A sky130_fd_sc_hd__inv_2
X_17693_ _17693_/A VGND VGND VPWR VPWR _17693_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15226__B1 _15208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19432_ _19431_/Y _19429_/X _19341_/X _19429_/X VGND VGND VPWR VPWR _23750_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13856_ _21386_/A _13852_/X _13524_/X _13852_/X VGND VGND VPWR VPWR _25261_/D sky130_fd_sc_hd__a2bb2o_4
X_16644_ _16182_/B _16643_/B VGND VGND VPWR VPWR _16644_/Y sky130_fd_sc_hd__nor2_4
X_12807_ _25385_/Q VGND VGND VPWR VPWR _12807_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19363_ _19362_/Y _19360_/X _19341_/X _19360_/X VGND VGND VPWR VPWR _19363_/X sky130_fd_sc_hd__a2bb2o_4
X_13787_ _14417_/A _14415_/A VGND VGND VPWR VPWR _14228_/A sky130_fd_sc_hd__or2_4
X_16575_ _16574_/Y _16572_/X _16315_/X _16572_/X VGND VGND VPWR VPWR _24543_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18314_ _21182_/A VGND VGND VPWR VPWR _18314_/X sky130_fd_sc_hd__buf_2
X_12738_ _12742_/A _12738_/B VGND VGND VPWR VPWR _12740_/B sky130_fd_sc_hd__or2_4
X_15526_ _15544_/A VGND VGND VPWR VPWR _15526_/X sky130_fd_sc_hd__buf_2
X_19294_ _21625_/B _19293_/X _16894_/X _19293_/X VGND VGND VPWR VPWR _23799_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21323__A1_N _17391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22138__A _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21042__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _14289_/X _20540_/B _15450_/Y _13950_/A _15453_/X VGND VGND VPWR VPWR _15457_/X
+ sky130_fd_sc_hd__a32o_4
X_18245_ _13828_/D VGND VGND VPWR VPWR _18245_/X sky130_fd_sc_hd__buf_2
X_12669_ _12636_/A _12669_/B _12668_/X VGND VGND VPWR VPWR _25429_/D sky130_fd_sc_hd__and3_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _25152_/Q VGND VGND VPWR VPWR _14408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15040__A _25023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21078__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15388_ _15388_/A _15314_/C VGND VGND VPWR VPWR _15389_/B sky130_fd_sc_hd__or2_4
X_18176_ _18037_/A _18174_/X _18175_/X VGND VGND VPWR VPWR _18176_/X sky130_fd_sc_hd__and3_4
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14339_ _14339_/A VGND VGND VPWR VPWR _14369_/A sky130_fd_sc_hd__buf_2
X_17127_ _17064_/A VGND VGND VPWR VPWR _17127_/X sky130_fd_sc_hd__buf_2
X_17058_ _17035_/Y _17057_/X VGND VGND VPWR VPWR _17068_/B sky130_fd_sc_hd__or2_4
XFILLER_171_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16009_ _16008_/Y _16006_/X _11755_/X _16006_/X VGND VGND VPWR VPWR _24751_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_HCLK clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__18651__B1 _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12279__B1 _12273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20971_ _20971_/A _13533_/A VGND VGND VPWR VPWR _24103_/D sky130_fd_sc_hd__nor2_4
XANTENNA__12839__A _25403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _22528_/X _22708_/X _22476_/A _22709_/X VGND VGND VPWR VPWR _22711_/A sky130_fd_sc_hd__o22a_4
X_23690_ _23690_/CLK _23690_/D VGND VGND VPWR VPWR _19605_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22641_ _22641_/A _21104_/B VGND VGND VPWR VPWR _22641_/X sky130_fd_sc_hd__or2_4
XANTENNA__14440__B2 _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25360_ _25358_/CLK _25360_/D HRESETn VGND VGND VPWR VPWR _25360_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17430__A _14423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22572_ _22289_/A _22571_/X _21550_/X _24731_/Q _21317_/X VGND VGND VPWR VPWR _22572_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16717__B1 _16537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24311_ _25543_/CLK _24311_/D HRESETn VGND VGND VPWR VPWR _17575_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_194_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21523_ _18278_/X _21518_/X _21520_/X _21522_/X VGND VGND VPWR VPWR _21524_/A sky130_fd_sc_hd__a211o_4
X_25291_ _25292_/CLK _25291_/D HRESETn VGND VGND VPWR VPWR _11685_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24242_ _24238_/CLK _24242_/D HRESETn VGND VGND VPWR VPWR _24242_/Q sky130_fd_sc_hd__dfrtp_4
X_21454_ _21711_/A _21447_/X _23321_/A _21453_/X VGND VGND VPWR VPWR _21454_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_108_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20405_ _20405_/A _21217_/A VGND VGND VPWR VPWR _20406_/A sky130_fd_sc_hd__or2_4
X_24173_ _24201_/CLK _18577_/X HRESETn VGND VGND VPWR VPWR _24173_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21385_ _21282_/X _21381_/X _21383_/Y _21384_/X VGND VGND VPWR VPWR _21385_/X sky130_fd_sc_hd__a211o_4
XFILLER_119_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_152_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _23631_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_162_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23124_ _22721_/B VGND VGND VPWR VPWR _23124_/X sky130_fd_sc_hd__buf_2
X_20336_ _20323_/Y VGND VGND VPWR VPWR _20336_/X sky130_fd_sc_hd__buf_2
XFILLER_1_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23055_ _23052_/X _23054_/X _22986_/X _24883_/Q _22784_/X VGND VGND VPWR VPWR _23056_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20267_ _13350_/B VGND VGND VPWR VPWR _20267_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22006_ _17900_/A _20356_/Y _22003_/X _22005_/X VGND VGND VPWR VPWR _22006_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20198_ _20193_/A VGND VGND VPWR VPWR _20198_/X sky130_fd_sc_hd__buf_2
XANTENNA__22511__A _15022_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11971_ _11712_/A _11968_/X _25507_/Q _11970_/X VGND VGND VPWR VPWR _25507_/D sky130_fd_sc_hd__o22a_4
X_23957_ _25137_/CLK _20591_/Y HRESETn VGND VGND VPWR VPWR _23957_/Q sky130_fd_sc_hd__dfrtp_4
X_13710_ _13710_/A VGND VGND VPWR VPWR _13710_/Y sky130_fd_sc_hd__inv_2
X_22908_ _22886_/X _22889_/X _22893_/Y _22907_/X VGND VGND VPWR VPWR HRDATA[18] sky130_fd_sc_hd__a211o_4
X_14690_ _21257_/A VGND VGND VPWR VPWR _22085_/A sky130_fd_sc_hd__buf_2
XFILLER_44_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23888_ _23459_/CLK _23888_/D VGND VGND VPWR VPWR _18125_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12468__B _13017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13641_ _19143_/A _13640_/X _19143_/A _13640_/X VGND VGND VPWR VPWR _13641_/X sky130_fd_sc_hd__a2bb2o_4
X_22839_ _21457_/X VGND VGND VPWR VPWR _22839_/X sky130_fd_sc_hd__buf_2
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23297__A3 _22145_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _16358_/Y _16359_/X _16070_/X _16359_/X VGND VGND VPWR VPWR _24623_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13572_ _13571_/Y _25102_/Q _13571_/Y _25102_/Q VGND VGND VPWR VPWR _13573_/D sky130_fd_sc_hd__a2bb2o_4
X_25558_ _25507_/CLK _25558_/D HRESETn VGND VGND VPWR VPWR _11712_/A sky130_fd_sc_hd__dfrtp_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15311_ _15311_/A VGND VGND VPWR VPWR _15423_/A sky130_fd_sc_hd__inv_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12523_ _24866_/Q VGND VGND VPWR VPWR _12523_/Y sky130_fd_sc_hd__inv_2
X_24509_ _24509_/CLK _16668_/X HRESETn VGND VGND VPWR VPWR _16666_/A sky130_fd_sc_hd__dfrtp_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16291_ _16291_/A VGND VGND VPWR VPWR _16291_/X sky130_fd_sc_hd__buf_2
XFILLER_188_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25489_ _25491_/CLK _12089_/X HRESETn VGND VGND VPWR VPWR _12087_/A sky130_fd_sc_hd__dfrtp_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15242_ _14969_/A _15241_/Y VGND VGND VPWR VPWR _15244_/B sky130_fd_sc_hd__or2_4
X_18030_ _15704_/X _18004_/X _18028_/X _24254_/Q _18029_/X VGND VGND VPWR VPWR _18030_/X
+ sky130_fd_sc_hd__o32a_4
X_12454_ _12208_/Y _12453_/X VGND VGND VPWR VPWR _12455_/C sky130_fd_sc_hd__nand2_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20268__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19122__B2 _19121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24855__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15173_ _15172_/X VGND VGND VPWR VPWR _15294_/A sky130_fd_sc_hd__buf_2
XFILLER_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15795__A _15934_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _12994_/A _12373_/Y _13004_/B _24829_/Q VGND VGND VPWR VPWR _12389_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14124_ _14124_/A _14124_/B _14110_/A VGND VGND VPWR VPWR _14125_/B sky130_fd_sc_hd__or3_4
X_19981_ _23558_/Q VGND VGND VPWR VPWR _19981_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15695__B1 _15694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14055_ _14054_/X VGND VGND VPWR VPWR _14055_/Y sky130_fd_sc_hd__inv_2
X_18932_ _21402_/B _18929_/X _16897_/X _18929_/X VGND VGND VPWR VPWR _23926_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13006_ _13006_/A _13006_/B _13006_/C VGND VGND VPWR VPWR _13052_/B sky130_fd_sc_hd__or3_4
XFILLER_239_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18863_ _24576_/Q _18683_/B _24576_/Q _18683_/B VGND VGND VPWR VPWR _18863_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11761__A1_N _11757_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17814_ _17770_/X _17780_/X _16952_/Y VGND VGND VPWR VPWR _17814_/X sky130_fd_sc_hd__o21a_4
XFILLER_223_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18794_ _18805_/A _18799_/B _18794_/C _18799_/C VGND VGND VPWR VPWR _18795_/A sky130_fd_sc_hd__or4_4
XANTENNA__15998__A1 _15797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17745_ _17710_/X _17898_/B _21834_/A VGND VGND VPWR VPWR _17909_/A sky130_fd_sc_hd__or3_4
X_14957_ _14956_/Y _16843_/A _14956_/Y _16843_/A VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13908_ _13908_/A VGND VGND VPWR VPWR _13963_/A sky130_fd_sc_hd__buf_2
X_17676_ _17522_/Y _17676_/B VGND VGND VPWR VPWR _17676_/X sky130_fd_sc_hd__or2_4
XANTENNA__12681__B1 _12657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16947__B1 _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14888_ _14888_/A VGND VGND VPWR VPWR _14888_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _19415_/A VGND VGND VPWR VPWR _19415_/X sky130_fd_sc_hd__buf_2
X_16627_ _16627_/A VGND VGND VPWR VPWR _16627_/Y sky130_fd_sc_hd__inv_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ _13589_/Y _13838_/X _11831_/X _13838_/X VGND VGND VPWR VPWR _25270_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19346_ _19346_/A _19346_/B _19346_/C VGND VGND VPWR VPWR _19346_/X sky130_fd_sc_hd__or3_4
X_16558_ _16558_/A VGND VGND VPWR VPWR _16558_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15509_ _15507_/Y _15508_/X HADDR[19] _15508_/X VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__a2bb2o_4
X_19277_ _23804_/Q VGND VGND VPWR VPWR _19277_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16489_ _16487_/Y _16483_/X _16402_/X _16488_/X VGND VGND VPWR VPWR _24576_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17372__B1 _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18228_ _18164_/A _23845_/Q VGND VGND VPWR VPWR _18230_/B sky130_fd_sc_hd__or2_4
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15201__C _15172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20259__B1 _19817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24596__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18159_ _18127_/A _18157_/X _18158_/X VGND VGND VPWR VPWR _18163_/B sky130_fd_sc_hd__and3_4
XANTENNA__24525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21170_ _21170_/A _21170_/B _21169_/X VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_225_0_HCLK clkbuf_7_112_0_HCLK/X VGND VGND VPWR VPWR _24334_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_172_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20121_ _23510_/Q VGND VGND VPWR VPWR _21418_/B sky130_fd_sc_hd__inv_2
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20052_ _20050_/Y _20051_/X _20007_/X _20051_/X VGND VGND VPWR VPWR _20052_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20431__B1 _20243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22971__A2 _22962_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24860_ _24872_/CLK _24860_/D HRESETn VGND VGND VPWR VPWR _24860_/Q sky130_fd_sc_hd__dfrtp_4
X_23811_ _23628_/CLK _23811_/D VGND VGND VPWR VPWR _23811_/Q sky130_fd_sc_hd__dfxtp_4
X_24791_ _24803_/CLK _15917_/X HRESETn VGND VGND VPWR VPWR _21432_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22184__B1 _25444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18927__B2 _18922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23742_ _23754_/CLK _19455_/X VGND VGND VPWR VPWR _18182_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _16662_/Y _20854_/A _20836_/A _20953_/Y VGND VGND VPWR VPWR _20954_/X sky130_fd_sc_hd__o22a_4
XFILLER_226_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16938__B1 _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23162__A _23162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23466_/CLK _23673_/D VGND VGND VPWR VPWR _13329_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _13670_/A VGND VGND VPWR VPWR _20885_/Y sky130_fd_sc_hd__inv_2
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15610__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25412_ _24476_/CLK _25412_/D HRESETn VGND VGND VPWR VPWR _25412_/Q sky130_fd_sc_hd__dfrtp_4
X_22624_ _22624_/A VGND VGND VPWR VPWR _22624_/Y sky130_fd_sc_hd__inv_2
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25343_ _25368_/CLK _13119_/X HRESETn VGND VGND VPWR VPWR _25343_/Q sky130_fd_sc_hd__dfrtp_4
X_22555_ _22528_/X _22551_/X _22431_/X _22554_/X VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21506_ _21468_/X _21506_/B VGND VGND VPWR VPWR _21507_/C sky130_fd_sc_hd__or2_4
X_25274_ _25103_/CLK _13833_/X HRESETn VGND VGND VPWR VPWR _25274_/Q sky130_fd_sc_hd__dfrtp_4
X_22486_ _21881_/X _22483_/X _22484_/X _24834_/Q _22485_/X VGND VGND VPWR VPWR _22486_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12304__A2_N _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24225_ _24238_/CLK _24225_/D HRESETn VGND VGND VPWR VPWR _24225_/Q sky130_fd_sc_hd__dfrtp_4
X_21437_ _21436_/X VGND VGND VPWR VPWR _22558_/A sky130_fd_sc_hd__buf_2
XFILLER_166_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16504__A _24569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _25171_/Q _12170_/B VGND VGND VPWR VPWR _12170_/X sky130_fd_sc_hd__or2_4
X_24156_ _23976_/CLK _24156_/D HRESETn VGND VGND VPWR VPWR _18681_/A sky130_fd_sc_hd__dfrtp_4
X_21368_ _14199_/B _21348_/B VGND VGND VPWR VPWR _21565_/A sky130_fd_sc_hd__or2_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18863__B1 _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23107_ _12781_/Y _22725_/X _22291_/B _12548_/Y _22862_/X VGND VGND VPWR VPWR _23107_/X
+ sky130_fd_sc_hd__o32a_4
X_20319_ _20319_/A VGND VGND VPWR VPWR _21200_/B sky130_fd_sc_hd__inv_2
X_24087_ _24339_/CLK _20539_/X HRESETn VGND VGND VPWR VPWR _24087_/Q sky130_fd_sc_hd__dfrtp_4
X_21299_ _21299_/A _15662_/Y _15673_/A _21109_/B VGND VGND VPWR VPWR _21597_/A sky130_fd_sc_hd__or4_4
X_23038_ _14980_/A _22851_/X _22108_/X _23037_/X VGND VGND VPWR VPWR _23038_/X sky130_fd_sc_hd__a211o_4
XFILLER_103_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15860_ _21173_/B VGND VGND VPWR VPWR _21592_/A sky130_fd_sc_hd__inv_2
X_14811_ _25056_/Q _14811_/B _14811_/C VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__or3_4
XFILLER_76_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15791_ _12059_/A _11721_/A _15791_/C _15791_/D VGND VGND VPWR VPWR _15792_/A sky130_fd_sc_hd__or4_4
X_24989_ _24989_/CLK _24989_/D HRESETn VGND VGND VPWR VPWR _24989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22714__A2 _22424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17530_ _25527_/Q _24298_/Q _11864_/Y _17529_/Y VGND VGND VPWR VPWR _17533_/C sky130_fd_sc_hd__o22a_4
XANTENNA__19550__A _16464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11954_ _20007_/A VGND VGND VPWR VPWR _19643_/A sky130_fd_sc_hd__buf_2
X_14742_ _14742_/A VGND VGND VPWR VPWR _14742_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19040__B1 _18969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12663__B1 _12662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14673_ _14672_/X VGND VGND VPWR VPWR _14674_/A sky130_fd_sc_hd__buf_2
X_17461_ _13211_/A _13410_/A VGND VGND VPWR VPWR _17461_/X sky130_fd_sc_hd__and2_4
X_11885_ _11885_/A _25516_/Q VGND VGND VPWR VPWR _11885_/X sky130_fd_sc_hd__and2_4
X_19200_ _19200_/A VGND VGND VPWR VPWR _19200_/Y sky130_fd_sc_hd__inv_2
X_13624_ _13613_/A VGND VGND VPWR VPWR _18102_/A sky130_fd_sc_hd__buf_2
X_16412_ HWDATA[20] VGND VGND VPWR VPWR _16412_/X sky130_fd_sc_hd__buf_2
XFILLER_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_234_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17392_ _17353_/A _17389_/B _17392_/C VGND VGND VPWR VPWR _24347_/D sky130_fd_sc_hd__and3_4
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ _19131_/A VGND VGND VPWR VPWR _19131_/X sky130_fd_sc_hd__buf_2
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13555_ _25272_/Q VGND VGND VPWR VPWR _13555_/Y sky130_fd_sc_hd__inv_2
X_16343_ _24629_/Q VGND VGND VPWR VPWR _16343_/Y sky130_fd_sc_hd__inv_2
X_12506_ _12505_/X VGND VGND VPWR VPWR _12506_/Y sky130_fd_sc_hd__inv_2
X_16274_ _16273_/Y _16269_/X _15995_/X _16269_/X VGND VGND VPWR VPWR _24654_/D sky130_fd_sc_hd__a2bb2o_4
X_19062_ _19060_/Y _19056_/X _19012_/X _19061_/X VGND VGND VPWR VPWR _23882_/D sky130_fd_sc_hd__a2bb2o_4
X_13486_ _13486_/A VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__buf_2
XFILLER_158_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15225_ _15252_/A _15223_/X _15224_/X VGND VGND VPWR VPWR _25034_/D sky130_fd_sc_hd__and3_4
X_18013_ _18013_/A VGND VGND VPWR VPWR _18200_/A sky130_fd_sc_hd__buf_2
XFILLER_172_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21320__A _21320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12437_ _12437_/A VGND VGND VPWR VPWR _12437_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16414__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15156_ _24605_/Q VGND VGND VPWR VPWR _15156_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12368_ _12997_/C _24840_/Q _12997_/C _24840_/Q VGND VGND VPWR VPWR _12369_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18854__B1 _16532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22650__B2 _22940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14107_ _14174_/A _14174_/B _14190_/A _14107_/D VGND VGND VPWR VPWR _14108_/B sky130_fd_sc_hd__or4_4
X_15087_ _25008_/Q VGND VGND VPWR VPWR _15340_/A sky130_fd_sc_hd__inv_2
X_19964_ _19964_/A VGND VGND VPWR VPWR _22353_/B sky130_fd_sc_hd__inv_2
XFILLER_180_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19725__A _19719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12299_ _12299_/A _12299_/B VGND VGND VPWR VPWR _12414_/A sky130_fd_sc_hd__or2_4
XFILLER_234_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14038_ _14013_/A _14013_/B _13999_/C _13999_/D VGND VGND VPWR VPWR _14039_/B sky130_fd_sc_hd__a211o_4
X_18915_ _19837_/A _20149_/B _18914_/X VGND VGND VPWR VPWR _18916_/A sky130_fd_sc_hd__or3_4
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19895_ _19895_/A VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_55_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24738_/CLK sky130_fd_sc_hd__clkbuf_1
X_18846_ _24561_/Q _24140_/Q _16524_/Y _18805_/A VGND VGND VPWR VPWR _18846_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18777_ _18772_/A _18772_/B _18740_/X _18773_/Y VGND VGND VPWR VPWR _18777_/X sky130_fd_sc_hd__a211o_4
X_15989_ _12190_/Y _15986_/X _15632_/X _15986_/X VGND VGND VPWR VPWR _15989_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15840__B1 _15629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17728_ _17723_/X _21675_/A _17723_/X _21675_/A VGND VGND VPWR VPWR _17743_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17659_ _17641_/A _17646_/D _17658_/X VGND VGND VPWR VPWR _24311_/D sky130_fd_sc_hd__and3_4
X_20670_ _14240_/Y _20622_/Y _20637_/A _20669_/X VGND VGND VPWR VPWR _20670_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23132__D _23131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24777__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19329_ _19328_/Y _19325_/X _19305_/X _19325_/X VGND VGND VPWR VPWR _19329_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11740__B _13786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21141__B2 _21353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18804__A _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24706__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22340_ _22339_/X VGND VGND VPWR VPWR _22340_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21230__A _21032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22271_ _22271_/A _22271_/B VGND VGND VPWR VPWR _22272_/C sky130_fd_sc_hd__or2_4
XFILLER_117_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16324__A _24636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24010_ _23980_/CLK _24010_/D HRESETn VGND VGND VPWR VPWR _24010_/Q sky130_fd_sc_hd__dfrtp_4
X_21222_ _24328_/Q _21222_/B VGND VGND VPWR VPWR _21222_/X sky130_fd_sc_hd__and2_4
XFILLER_145_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21153_ _21031_/X _21153_/B VGND VGND VPWR VPWR _21153_/Y sky130_fd_sc_hd__nor2_4
XFILLER_208_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20104_ _23515_/Q VGND VGND VPWR VPWR _20104_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21084_ _11747_/A VGND VGND VPWR VPWR _21085_/A sky130_fd_sc_hd__buf_2
XFILLER_247_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20035_ _20033_/Y _20029_/X _20034_/X _20016_/Y VGND VGND VPWR VPWR _20035_/X sky130_fd_sc_hd__a2bb2o_4
X_24912_ _24913_/CLK _24912_/D HRESETn VGND VGND VPWR VPWR _15611_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17281__C1 _17280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24843_ _25425_/CLK _15823_/X HRESETn VGND VGND VPWR VPWR _24843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15831__B1 _24838_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24774_ _24792_/CLK _24774_/D HRESETn VGND VGND VPWR VPWR _22982_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _20350_/Y _20343_/X VGND VGND VPWR VPWR _21986_/X sky130_fd_sc_hd__or2_4
XPHY_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _24217_/CLK _23725_/D VGND VGND VPWR VPWR _23725_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_82_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _20936_/Y _20933_/Y _13674_/X VGND VGND VPWR VPWR _20937_/X sky130_fd_sc_hd__o21a_4
XFILLER_27_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14398__B1 _13849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _24237_/Q VGND VGND VPWR VPWR _11670_/Y sky130_fd_sc_hd__inv_2
X_23656_ _23642_/CLK _23656_/D VGND VGND VPWR VPWR _13362_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _20867_/X VGND VGND VPWR VPWR _24054_/D sky130_fd_sc_hd__inv_2
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _21060_/A _22606_/X VGND VGND VPWR VPWR _22607_/Y sky130_fd_sc_hd__nand2_4
XFILLER_230_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21722__A1_N _12273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23587_ _23563_/CLK _23587_/D VGND VGND VPWR VPWR _19907_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17336__B1 _17288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ _15588_/Y _20716_/A _20724_/X _20798_/X VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__o22a_4
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13469_/A _13338_/X _13340_/C VGND VGND VPWR VPWR _13340_/X sky130_fd_sc_hd__and3_4
X_25326_ _25181_/CLK _13494_/X HRESETn VGND VGND VPWR VPWR _13493_/A sky130_fd_sc_hd__dfrtp_4
X_22538_ _22738_/A VGND VGND VPWR VPWR _23313_/B sky130_fd_sc_hd__buf_2
XFILLER_195_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22236__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15898__B1 _22755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13271_ _13271_/A VGND VGND VPWR VPWR _13411_/A sky130_fd_sc_hd__buf_2
X_25257_ _25204_/CLK _13874_/X HRESETn VGND VGND VPWR VPWR _13871_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22469_ _11695_/Y _21967_/A _13584_/Y _22523_/A VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__o22a_4
X_15010_ _15009_/X _23037_/A _15009_/X _23037_/A VGND VGND VPWR VPWR _15010_/X sky130_fd_sc_hd__a2bb2o_4
X_12222_ _25457_/Q VGND VGND VPWR VPWR _12222_/Y sky130_fd_sc_hd__inv_2
X_24208_ _23522_/CLK _18354_/Y HRESETn VGND VGND VPWR VPWR _13212_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25188_ _25188_/CLK _25188_/D HRESETn VGND VGND VPWR VPWR _25188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _25480_/Q _12152_/Y _25480_/Q _12152_/Y VGND VGND VPWR VPWR _12153_/X sky130_fd_sc_hd__a2bb2o_4
X_24139_ _25212_/CLK _24139_/D HRESETn VGND VGND VPWR VPWR _24139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12084_ _12072_/Y _12083_/X _11842_/X _12083_/X VGND VGND VPWR VPWR _12084_/X sky130_fd_sc_hd__a2bb2o_4
X_16961_ _16941_/X _16946_/X _16961_/C _16961_/D VGND VGND VPWR VPWR _16961_/X sky130_fd_sc_hd__or4_4
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18700_ _18700_/A _18700_/B VGND VGND VPWR VPWR _18733_/B sky130_fd_sc_hd__or2_4
X_15912_ _15875_/Y VGND VGND VPWR VPWR _15912_/X sky130_fd_sc_hd__buf_2
XFILLER_89_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17065__A _17393_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19680_ _19679_/Y _19676_/X _19656_/X _19676_/X VGND VGND VPWR VPWR _23667_/D sky130_fd_sc_hd__a2bb2o_4
X_16892_ _20122_/A VGND VGND VPWR VPWR _19810_/A sky130_fd_sc_hd__buf_2
XFILLER_238_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18631_ _16615_/A _24138_/Q _16615_/Y _18630_/Y VGND VGND VPWR VPWR _18631_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15843_ _12354_/Y _15842_/X _15636_/X _15842_/X VGND VGND VPWR VPWR _24830_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15822__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18562_ _18556_/X _18562_/B _18561_/X VGND VGND VPWR VPWR _24176_/D sky130_fd_sc_hd__and3_4
X_12986_ _12988_/A _12986_/B _12985_/Y VGND VGND VPWR VPWR _25374_/D sky130_fd_sc_hd__and3_4
X_15774_ _15751_/A VGND VGND VPWR VPWR _15774_/X sky130_fd_sc_hd__buf_2
XFILLER_206_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17513_ _25546_/Q _17579_/A _25552_/Q _17569_/B VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22163__A3 _22986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14725_ _22237_/A VGND VGND VPWR VPWR _14725_/X sky130_fd_sc_hd__buf_2
XANTENNA__21315__A _21332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11937_ _19993_/A VGND VGND VPWR VPWR _19629_/A sky130_fd_sc_hd__buf_2
X_18493_ _18493_/A VGND VGND VPWR VPWR _18828_/B sky130_fd_sc_hd__inv_2
XFILLER_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21371__A1 _14885_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11841__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17444_ _17443_/Y _17441_/X _16726_/X _17441_/X VGND VGND VPWR VPWR _17444_/X sky130_fd_sc_hd__a2bb2o_4
X_11868_ _11864_/Y _11857_/X _11867_/X _11857_/X VGND VGND VPWR VPWR _11868_/X sky130_fd_sc_hd__a2bb2o_4
X_14656_ _14656_/A VGND VGND VPWR VPWR _18130_/A sky130_fd_sc_hd__buf_2
XFILLER_21_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24870__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _13607_/A _13607_/B _25062_/Q _13606_/X VGND VGND VPWR VPWR _14679_/B sky130_fd_sc_hd__or4_4
XPHY_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17375_ _17378_/A _17378_/B VGND VGND VPWR VPWR _17375_/X sky130_fd_sc_hd__or2_4
XANTENNA__17327__B1 _17280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11799_ _25542_/Q VGND VGND VPWR VPWR _11799_/Y sky130_fd_sc_hd__inv_2
X_14587_ _25102_/Q _14586_/X _14584_/Y VGND VGND VPWR VPWR _25102_/D sky130_fd_sc_hd__o21a_4
XFILLER_41_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17428__A1_N _20680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19114_ _23862_/Q VGND VGND VPWR VPWR _21400_/B sky130_fd_sc_hd__inv_2
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16324_/Y _16320_/X _15967_/X _16325_/X VGND VGND VPWR VPWR _24636_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17878__A1 _16920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13538_ _13537_/X VGND VGND VPWR VPWR _13538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15138__A2_N _16432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15889__B1 _11790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19043_/Y _19044_/X _18975_/X _19044_/X VGND VGND VPWR VPWR _23887_/D sky130_fd_sc_hd__a2bb2o_4
X_13469_ _13469_/A _13467_/X _13469_/C VGND VGND VPWR VPWR _13470_/C sky130_fd_sc_hd__and3_4
X_16257_ _16264_/A VGND VGND VPWR VPWR _16257_/X sky130_fd_sc_hd__buf_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ _14996_/A VGND VGND VPWR VPWR _15208_/X sky130_fd_sc_hd__buf_2
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16188_ _14781_/A _16186_/Y _14772_/A _16186_/Y VGND VGND VPWR VPWR _16188_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22623__B2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20634__B1 _20680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15139_ _15139_/A VGND VGND VPWR VPWR _15139_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19947_ _22354_/B _19946_/X _19626_/X _19946_/X VGND VGND VPWR VPWR _23572_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19252__B1 _19184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19878_ _19878_/A VGND VGND VPWR VPWR _19878_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18829_ _18749_/A _18791_/B _18828_/X VGND VGND VPWR VPWR _24131_/D sky130_fd_sc_hd__and3_4
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11735__B _21135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15813__B1 _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21840_ _21833_/Y _21839_/X _21526_/X VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__o21a_4
XFILLER_243_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21771_ _21629_/A _21771_/B VGND VGND VPWR VPWR _21771_/X sky130_fd_sc_hd__or2_4
XANTENNA__21362__A1 SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16319__A _24638_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23510_ _23494_/CLK _23510_/D VGND VGND VPWR VPWR _23510_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20722_ _15631_/Y _20716_/X _20704_/X _20721_/Y VGND VGND VPWR VPWR _20722_/X sky130_fd_sc_hd__o22a_4
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24490_ _24493_/CLK _24490_/D HRESETn VGND VGND VPWR VPWR _16713_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_224_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23441_/CLK _23441_/D VGND VGND VPWR VPWR _23441_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20653_ _20653_/A _20651_/Y _20669_/C VGND VGND VPWR VPWR _20653_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_201_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14977__A2_N _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23372_ _23356_/X VGND VGND VPWR VPWR IRQ[16] sky130_fd_sc_hd__buf_2
XFILLER_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20584_ _20584_/A _18883_/B VGND VGND VPWR VPWR _20584_/Y sky130_fd_sc_hd__nand2_4
XFILLER_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25111_ _23970_/CLK _25111_/D HRESETn VGND VGND VPWR VPWR _25111_/Q sky130_fd_sc_hd__dfrtp_4
X_22323_ _14116_/A _17424_/A _20609_/A _22190_/B VGND VGND VPWR VPWR _22323_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25042_ _25043_/CLK _15190_/X HRESETn VGND VGND VPWR VPWR _15188_/A sky130_fd_sc_hd__dfrtp_4
X_22254_ _22265_/A _22252_/X _22253_/X VGND VGND VPWR VPWR _22254_/X sky130_fd_sc_hd__and3_4
XANTENNA__21895__A _21267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22614__B2 _22940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21205_ _21201_/X _21204_/X _22266_/A VGND VGND VPWR VPWR _21205_/X sky130_fd_sc_hd__o21a_4
XFILLER_191_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20625__B1 _20680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22185_ _21040_/Y _22184_/X VGND VGND VPWR VPWR _22185_/X sky130_fd_sc_hd__and2_4
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21136_ _21161_/A VGND VGND VPWR VPWR _21351_/A sky130_fd_sc_hd__inv_2
XFILLER_160_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21067_ _22694_/B VGND VGND VPWR VPWR _21067_/X sky130_fd_sc_hd__buf_2
XFILLER_247_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17316__C _17355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16057__B1 _11827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20018_ _22351_/B _20017_/X _19990_/X _20017_/X VGND VGND VPWR VPWR _23548_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12840_ _12839_/Y _23290_/A _12839_/Y _23290_/A VGND VGND VPWR VPWR _12840_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_246_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24826_ _24878_/CLK _15849_/X HRESETn VGND VGND VPWR VPWR _12353_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21135__A _21135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24699__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _12770_/Y _24790_/Q _12770_/Y _24790_/Q VGND VGND VPWR VPWR _12771_/X sky130_fd_sc_hd__a2bb2o_4
X_21969_ _21951_/X _21966_/X _21968_/X VGND VGND VPWR VPWR _21969_/X sky130_fd_sc_hd__a21o_4
X_24757_ _24757_/CLK _15992_/X HRESETn VGND VGND VPWR VPWR _24757_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_199_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11721_/Y VGND VGND VPWR VPWR _16190_/B sky130_fd_sc_hd__buf_2
X_14510_ _25116_/Q _14510_/B _14510_/C VGND VGND VPWR VPWR _14517_/A sky130_fd_sc_hd__or3_4
XFILLER_202_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24628__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _14890_/Y _15485_/X _15489_/X _15472_/A VGND VGND VPWR VPWR _15490_/X sky130_fd_sc_hd__a2bb2o_4
X_23708_ _23400_/CLK _23708_/D VGND VGND VPWR VPWR _22404_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_199_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24688_ _24712_/CLK _24688_/D HRESETn VGND VGND VPWR VPWR _21531_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_42_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _25142_/Q VGND VGND VPWR VPWR _14441_/Y sky130_fd_sc_hd__inv_2
X_23639_ _23631_/CLK _19757_/X VGND VGND VPWR VPWR _13401_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _14364_/X _14371_/X _12087_/A _14369_/X VGND VGND VPWR VPWR _14372_/X sky130_fd_sc_hd__o22a_4
X_17160_ _17139_/X _17160_/B _17160_/C VGND VGND VPWR VPWR _24383_/D sky130_fd_sc_hd__and3_4
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13323_ _13391_/A _13323_/B _13323_/C VGND VGND VPWR VPWR _13324_/C sky130_fd_sc_hd__or3_4
X_16111_ _16103_/X VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__buf_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25309_ _25309_/CLK _25309_/D HRESETn VGND VGND VPWR VPWR _25309_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17091_ _17088_/A _17088_/B VGND VGND VPWR VPWR _17091_/Y sky130_fd_sc_hd__nand2_4
XFILLER_171_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ _13451_/A VGND VGND VPWR VPWR _13254_/X sky130_fd_sc_hd__buf_2
X_16042_ _16042_/A VGND VGND VPWR VPWR _16042_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ _21083_/A VGND VGND VPWR VPWR _12205_/Y sky130_fd_sc_hd__inv_2
X_13185_ _13285_/A _13172_/X _13184_/X VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__or3_4
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19801_ _21899_/B _19797_/X _19800_/X _19797_/X VGND VGND VPWR VPWR _23625_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22413__B _21069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _12136_/A _12136_/B VGND VGND VPWR VPWR _12150_/A sky130_fd_sc_hd__and2_4
X_17993_ _18209_/A _23755_/Q VGND VGND VPWR VPWR _17996_/B sky130_fd_sc_hd__or2_4
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19732_ _13400_/B VGND VGND VPWR VPWR _19732_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12067_ _19594_/B VGND VGND VPWR VPWR _17448_/C sky130_fd_sc_hd__buf_2
X_16944_ _16132_/Y _16933_/A _22994_/A _17824_/A VGND VGND VPWR VPWR _16944_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19663_ _19662_/Y _19660_/X _19560_/X _19660_/X VGND VGND VPWR VPWR _23673_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19785__B2 _19765_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16875_ _16874_/X VGND VGND VPWR VPWR _16875_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23318__C1 _23317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18614_ _24141_/Q VGND VGND VPWR VPWR _18614_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_129_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _25062_/CLK sky130_fd_sc_hd__clkbuf_1
X_15826_ _15826_/A VGND VGND VPWR VPWR _15826_/X sky130_fd_sc_hd__buf_2
XFILLER_65_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19594_ _11731_/A _19594_/B _13786_/A _15670_/X VGND VGND VPWR VPWR _21161_/A sky130_fd_sc_hd__or4_4
XFILLER_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23244__B _23303_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ _18540_/A _18548_/B VGND VGND VPWR VPWR _18546_/C sky130_fd_sc_hd__nand2_4
X_15757_ _15737_/X _15751_/X _15756_/X _24873_/Q _15749_/X VGND VGND VPWR VPWR _15757_/X
+ sky130_fd_sc_hd__a32o_4
X_12969_ _12969_/A _12969_/B VGND VGND VPWR VPWR _12969_/X sky130_fd_sc_hd__or2_4
XFILLER_80_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17548__B1 _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _14723_/A VGND VGND VPWR VPWR _21262_/A sky130_fd_sc_hd__inv_2
X_18476_ _18476_/A _18476_/B _18418_/Y _18400_/Y VGND VGND VPWR VPWR _18476_/X sky130_fd_sc_hd__or4_4
X_15688_ _24894_/Q VGND VGND VPWR VPWR _15691_/C sky130_fd_sc_hd__inv_2
XANTENNA__16220__B1 _15960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15023__B2 _15022_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17427_ _14420_/A VGND VGND VPWR VPWR _17427_/X sky130_fd_sc_hd__buf_2
XANTENNA__23260__A _16201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14639_ _14639_/A _14639_/B VGND VGND VPWR VPWR _14639_/Y sky130_fd_sc_hd__nor2_4
XFILLER_220_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17358_ _17198_/X _17378_/A _17358_/C _17380_/A VGND VGND VPWR VPWR _17364_/C sky130_fd_sc_hd__or4_4
XFILLER_146_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16309_ HWDATA[25] VGND VGND VPWR VPWR _16309_/X sky130_fd_sc_hd__buf_2
X_17289_ _17243_/X _17277_/X _17288_/X _17284_/Y VGND VGND VPWR VPWR _17289_/X sky130_fd_sc_hd__a211o_4
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19028_ _19143_/A _19028_/B _19028_/C VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__or3_4
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25306__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11746__A _22575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23990_ _23991_/CLK _20641_/Y HRESETn VGND VGND VPWR VPWR _17399_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16039__B1 _15970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_25_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22941_ _22941_/A VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__buf_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_88_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_88_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18529__A _18515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22780__B1 _24841_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17433__A _14427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22872_ _22157_/C VGND VGND VPWR VPWR _22872_/X sky130_fd_sc_hd__buf_2
X_21823_ _22029_/A _21821_/X _21822_/X VGND VGND VPWR VPWR _21823_/X sky130_fd_sc_hd__and3_4
X_24611_ _24613_/CLK _24611_/D HRESETn VGND VGND VPWR VPWR _24611_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24792__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17539__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24721__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24542_ _24542_/CLK _24542_/D HRESETn VGND VGND VPWR VPWR _16576_/A sky130_fd_sc_hd__dfrtp_4
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21754_ _22459_/A _21751_/X _22462_/A _21753_/X VGND VGND VPWR VPWR _21755_/B sky130_fd_sc_hd__o22a_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21886__A2 _21436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16211__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20705_ _13130_/Y _13132_/B _13134_/B VGND VGND VPWR VPWR _20705_/X sky130_fd_sc_hd__o21a_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24473_ _24473_/CLK _24473_/D HRESETn VGND VGND VPWR VPWR _23037_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23088__A1 _16571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21685_ _21209_/A VGND VGND VPWR VPWR _21685_/X sky130_fd_sc_hd__buf_2
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23424_ _23400_/CLK _23424_/D VGND VGND VPWR VPWR _23424_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20636_ _14816_/A VGND VGND VPWR VPWR _20637_/A sky130_fd_sc_hd__buf_2
XANTENNA__22835__A1 _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23355_ _25279_/Q _21982_/X _23353_/Y _23354_/Y VGND VGND VPWR VPWR _23356_/B sky130_fd_sc_hd__a211o_4
XFILLER_166_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20567_ _20567_/A _20566_/Y _20556_/X VGND VGND VPWR VPWR _20567_/X sky130_fd_sc_hd__and3_4
XFILLER_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22306_ _22306_/A VGND VGND VPWR VPWR _22306_/X sky130_fd_sc_hd__buf_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23286_ _23263_/X _23267_/X _23286_/C _23285_/X VGND VGND VPWR VPWR HRDATA[29] sky130_fd_sc_hd__or4_4
X_20498_ _20493_/X _20497_/X VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__or2_4
XANTENNA__16514__A1_N _16512_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22599__B1 _22431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25025_ _25023_/CLK _15254_/Y HRESETn VGND VGND VPWR VPWR _14956_/A sky130_fd_sc_hd__dfrtp_4
X_22237_ _22237_/A _22229_/X _22236_/X VGND VGND VPWR VPWR _22237_/X sky130_fd_sc_hd__and3_4
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19464__B1 _19418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22168_ _24591_/Q _22945_/A VGND VGND VPWR VPWR _22171_/B sky130_fd_sc_hd__or2_4
XFILLER_121_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21119_ _13131_/B VGND VGND VPWR VPWR _21119_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23012__A1 _16578_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ _14990_/A VGND VGND VPWR VPWR _14990_/X sky130_fd_sc_hd__buf_2
X_22099_ _21785_/X _22098_/X _21277_/A VGND VGND VPWR VPWR _22099_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_219_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13941_ _24979_/Q VGND VGND VPWR VPWR _13941_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24809__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _16654_/X VGND VGND VPWR VPWR _16660_/X sky130_fd_sc_hd__buf_2
X_13872_ _13872_/A VGND VGND VPWR VPWR _13872_/X sky130_fd_sc_hd__buf_2
XFILLER_219_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15611_ _15611_/A VGND VGND VPWR VPWR _15611_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23315__A2 _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12823_ _12912_/A _22755_/A _12912_/A _22755_/A VGND VGND VPWR VPWR _12823_/X sky130_fd_sc_hd__a2bb2o_4
X_24809_ _24812_/CLK _24809_/D HRESETn VGND VGND VPWR VPWR _22913_/A sky130_fd_sc_hd__dfrtp_4
X_16591_ _16623_/A VGND VGND VPWR VPWR _16618_/A sky130_fd_sc_hd__buf_2
XANTENNA__21326__A1 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18330_ _20079_/A VGND VGND VPWR VPWR _18938_/A sky130_fd_sc_hd__buf_2
XFILLER_203_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _21140_/A VGND VGND VPWR VPWR _16462_/C sky130_fd_sc_hd__inv_2
X_12754_ _12869_/A _24821_/Q _12869_/A _24821_/Q VGND VGND VPWR VPWR _12760_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11705_/A VGND VGND VPWR VPWR _11705_/Y sky130_fd_sc_hd__inv_2
X_18261_ _18245_/X _18247_/X _15775_/X _24235_/Q _18248_/X VGND VGND VPWR VPWR _24235_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12619_/A _12619_/B _12618_/B _12685_/D VGND VGND VPWR VPWR _12691_/B sky130_fd_sc_hd__or4_4
X_15473_ _15470_/Y _15472_/X _14420_/X _15472_/X VGND VGND VPWR VPWR _15473_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17212_/A VGND VGND VPWR VPWR _17330_/A sky130_fd_sc_hd__inv_2
XANTENNA__22408__B _21656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _14137_/Y _14418_/X _14423_/X _14418_/X VGND VGND VPWR VPWR _14424_/X sky130_fd_sc_hd__a2bb2o_4
X_18192_ _18060_/A _18192_/B VGND VGND VPWR VPWR _18194_/B sky130_fd_sc_hd__or2_4
XANTENNA__21312__B _21312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _16992_/Y _17142_/X VGND VGND VPWR VPWR _17143_/X sky130_fd_sc_hd__or2_4
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _14349_/A _14359_/B _14334_/X VGND VGND VPWR VPWR _14355_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18902__A _14388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14207__A _14816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13306_ _13306_/A VGND VGND VPWR VPWR _13456_/A sky130_fd_sc_hd__buf_2
X_14286_ _23979_/Q VGND VGND VPWR VPWR _14286_/Y sky130_fd_sc_hd__inv_2
X_17074_ _17074_/A _17345_/A VGND VGND VPWR VPWR _17074_/X sky130_fd_sc_hd__and2_4
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18650__A1_N _16601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13237_ _13282_/A _23523_/Q VGND VGND VPWR VPWR _13237_/X sky130_fd_sc_hd__or2_4
X_16025_ _16023_/Y _16019_/X _15957_/X _16024_/X VGND VGND VPWR VPWR _16025_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19455__B1 _19454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16422__A _16390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13168_ _13192_/A _23676_/Q VGND VGND VPWR VPWR _13168_/X sky130_fd_sc_hd__or2_4
X_12119_ _12118_/Y _12116_/X _11847_/X _12116_/X VGND VGND VPWR VPWR _25480_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19733__A _19719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ _13002_/D _13102_/B VGND VGND VPWR VPWR _13100_/C sky130_fd_sc_hd__nand2_4
X_17976_ _13613_/B VGND VGND VPWR VPWR _17977_/A sky130_fd_sc_hd__buf_2
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21553__A1_N _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19715_ _13458_/B VGND VGND VPWR VPWR _19715_/Y sky130_fd_sc_hd__inv_2
X_16927_ _17871_/A VGND VGND VPWR VPWR _17861_/A sky130_fd_sc_hd__inv_2
XFILLER_226_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18349__A _17461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19646_ _19646_/A VGND VGND VPWR VPWR _19646_/X sky130_fd_sc_hd__buf_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16858_ _16856_/Y _16853_/X _16791_/X _16857_/X VGND VGND VPWR VPWR _24423_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16441__B1 _16066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15809_ _12337_/Y _15808_/X _11758_/X _15808_/X VGND VGND VPWR VPWR _24854_/D sky130_fd_sc_hd__a2bb2o_4
X_19577_ _23699_/Q VGND VGND VPWR VPWR _22247_/B sky130_fd_sc_hd__inv_2
X_16789_ _15000_/Y _16787_/X _16537_/X _16787_/X VGND VGND VPWR VPWR _24456_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22514__B1 _21591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18528_ _18493_/A VGND VGND VPWR VPWR _18550_/A sky130_fd_sc_hd__buf_2
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21503__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18459_ _18733_/C VGND VGND VPWR VPWR _18710_/A sky130_fd_sc_hd__buf_2
XFILLER_178_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18084__A _18008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21470_ _21815_/A _21467_/X _21469_/X VGND VGND VPWR VPWR _21470_/X sky130_fd_sc_hd__and3_4
X_20421_ _23395_/Q _20420_/Y _20994_/A _20419_/X VGND VGND VPWR VPWR _20421_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16943__A2_N _17751_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23140_ _15583_/Y _23140_/B VGND VGND VPWR VPWR _23140_/X sky130_fd_sc_hd__and2_4
X_20352_ _20352_/A VGND VGND VPWR VPWR _20352_/X sky130_fd_sc_hd__buf_2
XFILLER_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23071_ _22801_/X _23069_/X _22804_/X _23070_/X VGND VGND VPWR VPWR _23072_/B sky130_fd_sc_hd__o22a_4
X_20283_ _23450_/Q VGND VGND VPWR VPWR _22085_/B sky130_fd_sc_hd__inv_2
XANTENNA__16332__A _16290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22022_ _22034_/A _22022_/B VGND VGND VPWR VPWR _22025_/B sky130_fd_sc_hd__or2_4
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19643__A _19643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23973_ _23973_/CLK _23973_/D HRESETn VGND VGND VPWR VPWR _21020_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13494__B1 _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24902__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22924_ _22204_/A VGND VGND VPWR VPWR _22924_/X sky130_fd_sc_hd__buf_2
XFILLER_216_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_112_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _24825_/CLK sky130_fd_sc_hd__clkbuf_1
X_22855_ _14950_/A _22851_/X _22852_/X _22854_/X VGND VGND VPWR VPWR _22855_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22505__B1 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_175_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _24111_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21806_ _21668_/A _21806_/B VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__or2_4
XFILLER_225_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22786_ _23056_/A _22786_/B VGND VGND VPWR VPWR _22786_/X sky130_fd_sc_hd__and2_4
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21737_ _14225_/Y _14202_/X _14242_/Y _21356_/X VGND VGND VPWR VPWR _21738_/A sky130_fd_sc_hd__o22a_4
X_24525_ _24528_/CLK _24525_/D HRESETn VGND VGND VPWR VPWR _16620_/A sky130_fd_sc_hd__dfrtp_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16735__B2 _16734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12470_ _12469_/X VGND VGND VPWR VPWR _12470_/Y sky130_fd_sc_hd__inv_2
X_21668_ _21668_/A _19894_/Y VGND VGND VPWR VPWR _21670_/B sky130_fd_sc_hd__or2_4
X_24456_ _24430_/CLK _24456_/D HRESETn VGND VGND VPWR VPWR _24456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20619_ _20480_/X _20513_/X VGND VGND VPWR VPWR _23972_/D sky130_fd_sc_hd__and2_4
X_23407_ _23407_/CLK _23407_/D VGND VGND VPWR VPWR _23407_/Q sky130_fd_sc_hd__dfxtp_4
X_24387_ _24383_/CLK _17150_/X HRESETn VGND VGND VPWR VPWR _24387_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19685__B1 _19560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21599_ _15650_/X VGND VGND VPWR VPWR _21606_/A sky130_fd_sc_hd__buf_2
XFILLER_137_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16453__A1_N _15134_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ _14134_/X _14139_/X _25229_/Q _14134_/X VGND VGND VPWR VPWR _14140_/X sky130_fd_sc_hd__a2bb2o_4
X_23338_ _22535_/B _23338_/B VGND VGND VPWR VPWR _23338_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17696__C1 _17611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14071_ _13985_/X VGND VGND VPWR VPWR _20470_/B sky130_fd_sc_hd__inv_2
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23269_ _12225_/Y _22507_/X _23268_/X VGND VGND VPWR VPWR _23269_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12770__A _21035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ _13022_/A VGND VGND VPWR VPWR _13022_/Y sky130_fd_sc_hd__inv_2
X_25008_ _25002_/CLK _15341_/X HRESETn VGND VGND VPWR VPWR _25008_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17830_ _16923_/Y _17834_/B _17829_/Y VGND VGND VPWR VPWR _17830_/X sky130_fd_sc_hd__o21a_4
XFILLER_126_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17761_ _16920_/Y _16901_/Y _17761_/C _17761_/D VGND VGND VPWR VPWR _17761_/X sky130_fd_sc_hd__or4_4
X_14973_ _25035_/Q VGND VGND VPWR VPWR _14973_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14697__A _21263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19500_ _23725_/Q VGND VGND VPWR VPWR _21190_/B sky130_fd_sc_hd__inv_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16712_ _16711_/Y _16709_/X _16530_/X _16709_/X VGND VGND VPWR VPWR _16712_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24643__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _24980_/Q _13924_/B _13924_/C _13924_/D VGND VGND VPWR VPWR _13924_/X sky130_fd_sc_hd__or4_4
X_17692_ _17676_/B _17690_/Y _17702_/C VGND VGND VPWR VPWR _17692_/X sky130_fd_sc_hd__and3_4
XANTENNA__21307__B _21307_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_71_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19431_ _18181_/B VGND VGND VPWR VPWR _19431_/Y sky130_fd_sc_hd__inv_2
X_16643_ _16643_/A _16643_/B VGND VGND VPWR VPWR _16643_/X sky130_fd_sc_hd__or2_4
XFILLER_207_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13855_ _25261_/Q VGND VGND VPWR VPWR _21386_/A sky130_fd_sc_hd__inv_2
X_12806_ _12853_/A _12804_/Y _25378_/Q _12805_/Y VGND VGND VPWR VPWR _12806_/X sky130_fd_sc_hd__a2bb2o_4
X_19362_ _18192_/B VGND VGND VPWR VPWR _19362_/Y sky130_fd_sc_hd__inv_2
X_16574_ _16574_/A VGND VGND VPWR VPWR _16574_/Y sky130_fd_sc_hd__inv_2
X_13786_ _13786_/A VGND VGND VPWR VPWR _14415_/A sky130_fd_sc_hd__buf_2
XFILLER_15_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18313_ _24217_/Q VGND VGND VPWR VPWR _21182_/A sky130_fd_sc_hd__inv_2
X_15525_ _15499_/A VGND VGND VPWR VPWR _15544_/A sky130_fd_sc_hd__buf_2
X_12737_ _12737_/A _12737_/B VGND VGND VPWR VPWR _12738_/B sky130_fd_sc_hd__or2_4
X_19293_ _19280_/Y VGND VGND VPWR VPWR _19293_/X sky130_fd_sc_hd__buf_2
XFILLER_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16417__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18244_ _22745_/A _18243_/X _15752_/X _18243_/X VGND VGND VPWR VPWR _24246_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15456_ _13950_/A _15446_/X _15455_/X _13951_/B _15453_/X VGND VGND VPWR VPWR _15456_/X
+ sky130_fd_sc_hd__a32o_4
X_12668_ _25429_/Q _12671_/B VGND VGND VPWR VPWR _12668_/X sky130_fd_sc_hd__or2_4
XFILLER_31_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _14406_/Y _14403_/X _14248_/X _14392_/X VGND VGND VPWR VPWR _25153_/D sky130_fd_sc_hd__a2bb2o_4
X_18175_ _18036_/A _18175_/B VGND VGND VPWR VPWR _18175_/X sky130_fd_sc_hd__or2_4
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19728__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15387_ _15387_/A VGND VGND VPWR VPWR _15393_/A sky130_fd_sc_hd__buf_2
X_12599_ _12599_/A VGND VGND VPWR VPWR _12599_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17126_ _17126_/A VGND VGND VPWR VPWR _24392_/D sky130_fd_sc_hd__inv_2
X_14338_ _14338_/A _14359_/A VGND VGND VPWR VPWR _14339_/A sky130_fd_sc_hd__or2_4
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17057_ _17057_/A _17057_/B _17057_/C _17057_/D VGND VGND VPWR VPWR _17057_/X sky130_fd_sc_hd__or4_4
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17248__A _17305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14269_ _14263_/Y _14268_/X _13844_/X _14268_/X VGND VGND VPWR VPWR _14269_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16152__A _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16008_ _16008_/A VGND VGND VPWR VPWR _16008_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15600__A1_N _22934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22601__B _16382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17959_ _17944_/A _20232_/A VGND VGND VPWR VPWR _17960_/C sky130_fd_sc_hd__or2_4
XANTENNA__12279__B2 _21715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18079__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20970_ _24247_/Q _14628_/Y _15923_/B _13548_/A _15694_/X VGND VGND VPWR VPWR _20970_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_54_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21217__B _21351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25137__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19629_ _19629_/A VGND VGND VPWR VPWR _19629_/X sky130_fd_sc_hd__buf_2
XFILLER_54_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22640_ _22754_/A _22640_/B _22639_/X VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__and3_4
XANTENNA__13016__A _13049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_248_0_HCLK clkbuf_8_249_0_HCLK/A VGND VGND VPWR VPWR _24000_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23160__B1 _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22571_ _16348_/A _22610_/B VGND VGND VPWR VPWR _22571_/X sky130_fd_sc_hd__or2_4
XFILLER_222_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12855__A _12855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16327__A _24635_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21710__B2 _22530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21522_ _11661_/A _22062_/A VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__and2_4
X_24310_ _25520_/CLK _17661_/Y HRESETn VGND VGND VPWR VPWR _24310_/Q sky130_fd_sc_hd__dfrtp_4
X_25290_ _25292_/CLK _25290_/D HRESETn VGND VGND VPWR VPWR _11665_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16882__A2_N _16877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24241_ _24240_/CLK _24241_/D HRESETn VGND VGND VPWR VPWR _24241_/Q sky130_fd_sc_hd__dfrtp_4
X_21453_ _21307_/B _21451_/X _21314_/X _12353_/A _22531_/B VGND VGND VPWR VPWR _21453_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20404_ _21382_/B VGND VGND VPWR VPWR _20404_/X sky130_fd_sc_hd__buf_2
X_24172_ _24169_/CLK _24172_/D HRESETn VGND VGND VPWR VPWR _18423_/A sky130_fd_sc_hd__dfrtp_4
X_21384_ _13815_/Y _21384_/B VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__and2_4
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23123_ _21321_/X VGND VGND VPWR VPWR _23123_/X sky130_fd_sc_hd__buf_2
X_20335_ _20335_/A VGND VGND VPWR VPWR _21683_/B sky130_fd_sc_hd__inv_2
XANTENNA__19419__B1 _19418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23054_ _23054_/A _23119_/B VGND VGND VPWR VPWR _23054_/X sky130_fd_sc_hd__or2_4
XFILLER_150_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20266_ _20265_/Y _20263_/X _20243_/X _20263_/X VGND VGND VPWR VPWR _20266_/X sky130_fd_sc_hd__a2bb2o_4
X_22005_ _22005_/A _20360_/Y _22004_/X VGND VGND VPWR VPWR _22005_/X sky130_fd_sc_hd__and3_4
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20197_ _23482_/Q VGND VGND VPWR VPWR _20197_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22511__B _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11970_ _25506_/Q _25505_/Q _11970_/C _11970_/D VGND VGND VPWR VPWR _11970_/X sky130_fd_sc_hd__and4_4
X_23956_ _25137_/CLK _23956_/D HRESETn VGND VGND VPWR VPWR _20584_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_217_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_58_0_HCLK clkbuf_6_58_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20201__B2 _20198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22907_ _23020_/A _22895_/Y _22900_/X _22907_/D VGND VGND VPWR VPWR _22907_/X sky130_fd_sc_hd__or4_4
XFILLER_232_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23887_ _23889_/CLK _23887_/D VGND VGND VPWR VPWR _18157_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16956__B2 _24293_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13640_ _18089_/A _13615_/A _13639_/X _13615_/Y VGND VGND VPWR VPWR _13640_/X sky130_fd_sc_hd__o22a_4
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22838_ _22732_/A VGND VGND VPWR VPWR _23280_/A sky130_fd_sc_hd__buf_2
XFILLER_112_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _25274_/Q VGND VGND VPWR VPWR _13571_/Y sky130_fd_sc_hd__inv_2
X_25557_ _25507_/CLK _25557_/D HRESETn VGND VGND VPWR VPWR _11656_/A sky130_fd_sc_hd__dfrtp_4
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ _21440_/X _22764_/X _21844_/X _22768_/Y VGND VGND VPWR VPWR _22769_/X sky130_fd_sc_hd__a211o_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12765__A _25399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21701__B2 _21656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15310_ _15310_/A _15424_/A _15082_/Y _15407_/A VGND VGND VPWR VPWR _15310_/X sky130_fd_sc_hd__or4_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12521_/Y _24891_/Q _12521_/Y _24891_/Q VGND VGND VPWR VPWR _12522_/X sky130_fd_sc_hd__a2bb2o_4
X_24508_ _24073_/CLK _16670_/X HRESETn VGND VGND VPWR VPWR _16669_/A sky130_fd_sc_hd__dfrtp_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ _16290_/A VGND VGND VPWR VPWR _16291_/A sky130_fd_sc_hd__buf_2
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25488_ _25488_/CLK _12091_/X HRESETn VGND VGND VPWR VPWR _12090_/A sky130_fd_sc_hd__dfrtp_4
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _15240_/X VGND VGND VPWR VPWR _15241_/Y sky130_fd_sc_hd__inv_2
X_12453_ _12255_/Y _12453_/B VGND VGND VPWR VPWR _12453_/X sky130_fd_sc_hd__or2_4
X_24439_ _24437_/CLK _24439_/D HRESETn VGND VGND VPWR VPWR _14978_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19548__A _19548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12384_ _13011_/A _24855_/Q _13011_/A _24855_/Q VGND VGND VPWR VPWR _12384_/X sky130_fd_sc_hd__a2bb2o_4
X_15172_ _15172_/A _15171_/X VGND VGND VPWR VPWR _15172_/X sky130_fd_sc_hd__or2_4
XFILLER_126_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14123_ _14108_/C _14122_/X _25221_/Q VGND VGND VPWR VPWR _14124_/B sky130_fd_sc_hd__or3_4
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17068__A _17074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19980_ _21675_/B _19979_/X _19643_/X _19979_/X VGND VGND VPWR VPWR _23559_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18931_ _18931_/A VGND VGND VPWR VPWR _21402_/B sky130_fd_sc_hd__inv_2
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24895__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14054_ _14042_/X _14053_/X _14054_/C _14001_/X VGND VGND VPWR VPWR _14054_/X sky130_fd_sc_hd__or4_4
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22702__A _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13005_ _13005_/A _13002_/X _13004_/X VGND VGND VPWR VPWR _13006_/C sky130_fd_sc_hd__or3_4
XANTENNA__24824__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ _16532_/A _18810_/A _16519_/Y _18604_/X VGND VGND VPWR VPWR _18862_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19830__B1 _19734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17813_ _17748_/X _17803_/X _17813_/C VGND VGND VPWR VPWR _24286_/D sky130_fd_sc_hd__and3_4
X_18793_ _18630_/Y _18810_/A _18809_/A _18809_/B VGND VGND VPWR VPWR _18799_/C sky130_fd_sc_hd__or4_4
XFILLER_239_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15998__A2 _15895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11844__A _25531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17744_ _17743_/X VGND VGND VPWR VPWR _17744_/Y sky130_fd_sc_hd__inv_2
X_14956_ _14956_/A VGND VGND VPWR VPWR _14956_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13907_ _13927_/B VGND VGND VPWR VPWR _13907_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17675_ _17504_/Y _17674_/X VGND VGND VPWR VPWR _17676_/B sky130_fd_sc_hd__or2_4
XFILLER_223_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14887_ _14885_/Y _14819_/X _14844_/X _14886_/Y VGND VGND VPWR VPWR _14888_/A sky130_fd_sc_hd__o22a_4
XFILLER_208_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19414_ _19413_/X VGND VGND VPWR VPWR _19415_/A sky130_fd_sc_hd__inv_2
X_16626_ _16625_/Y _16623_/X _16368_/X _16623_/X VGND VGND VPWR VPWR _16626_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13838_ _13838_/A VGND VGND VPWR VPWR _13838_/X sky130_fd_sc_hd__buf_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16975__A1_N _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19345_ _17943_/B VGND VGND VPWR VPWR _19345_/Y sky130_fd_sc_hd__inv_2
X_16557_ _16556_/Y _16554_/X _16294_/X _16554_/X VGND VGND VPWR VPWR _24550_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_1_0_HCLK clkbuf_7_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13769_ _25284_/Q _13767_/B _13768_/Y VGND VGND VPWR VPWR _13769_/X sky130_fd_sc_hd__o21a_4
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_15_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _24295_/CLK sky130_fd_sc_hd__clkbuf_1
X_15508_ _15503_/A VGND VGND VPWR VPWR _15508_/X sky130_fd_sc_hd__buf_2
X_19276_ _21243_/B _19271_/X _18934_/X _19258_/Y VGND VGND VPWR VPWR _23805_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16488_ _16495_/A VGND VGND VPWR VPWR _16488_/X sky130_fd_sc_hd__buf_2
XANTENNA__17372__A1 _17364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_78_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24767_/CLK sky130_fd_sc_hd__clkbuf_1
X_18227_ _18227_/A _18227_/B _18227_/C VGND VGND VPWR VPWR _18227_/X sky130_fd_sc_hd__or3_4
X_15439_ _24005_/Q _23979_/Q _14257_/D _15444_/A VGND VGND VPWR VPWR _15439_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18158_ _18158_/A _19067_/A VGND VGND VPWR VPWR _18158_/X sky130_fd_sc_hd__or2_4
XFILLER_190_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17109_ _17042_/D _17101_/B VGND VGND VPWR VPWR _17110_/B sky130_fd_sc_hd__or2_4
X_18089_ _18089_/A VGND VGND VPWR VPWR _18107_/A sky130_fd_sc_hd__buf_2
X_20120_ _20117_/Y _20118_/X _20119_/X _20118_/X VGND VGND VPWR VPWR _23511_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24565__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20051_ _20038_/Y VGND VGND VPWR VPWR _20051_/X sky130_fd_sc_hd__buf_2
XANTENNA__16610__A _16618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17425__B _14232_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23810_ _23628_/CLK _23810_/D VGND VGND VPWR VPWR _19263_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_100_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16650__A3 HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24790_ _24825_/CLK _15918_/X HRESETn VGND VGND VPWR VPWR _24790_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12121__B1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22184__B2 _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _24074_/Q _20949_/X _20952_/Y VGND VGND VPWR VPWR _20953_/Y sky130_fd_sc_hd__a21oi_4
X_23741_ _23754_/CLK _23741_/D VGND VGND VPWR VPWR _18214_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20878_/X _20880_/Y _24494_/Q _20883_/X VGND VGND VPWR VPWR _24057_/D sky130_fd_sc_hd__a2bb2o_4
X_23672_ _23466_/CLK _23672_/D VGND VGND VPWR VPWR _13365_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_198_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23133__B1 _17752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25411_ _25410_/CLK _12734_/X HRESETn VGND VGND VPWR VPWR _25411_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _22607_/Y _22612_/Y _22620_/Y _21455_/X _22622_/X VGND VGND VPWR VPWR _22624_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22554_ _17359_/C _22677_/B _22553_/Y VGND VGND VPWR VPWR _22554_/X sky130_fd_sc_hd__o21a_4
X_25342_ _25368_/CLK _13121_/X HRESETn VGND VGND VPWR VPWR _12342_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21898__A _21263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21505_ _21668_/A _21505_/B VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__or2_4
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22485_ _11747_/A VGND VGND VPWR VPWR _22485_/X sky130_fd_sc_hd__buf_2
X_25273_ _25103_/CLK _13835_/X HRESETn VGND VGND VPWR VPWR _13578_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21447__B1 _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21436_ _22578_/B VGND VGND VPWR VPWR _21436_/X sky130_fd_sc_hd__buf_2
X_24224_ _24295_/CLK _18291_/X HRESETn VGND VGND VPWR VPWR _24224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24155_ _23976_/CLK _18742_/Y HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_238_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21367_ _21366_/X VGND VGND VPWR VPWR _21367_/Y sky130_fd_sc_hd__inv_2
X_20318_ _21469_/B _20315_/X _20010_/X _20315_/X VGND VGND VPWR VPWR _20318_/X sky130_fd_sc_hd__a2bb2o_4
X_23106_ _23106_/A _23105_/X VGND VGND VPWR VPWR _23106_/Y sky130_fd_sc_hd__nor2_4
X_24086_ _24339_/CLK _20538_/X HRESETn VGND VGND VPWR VPWR _24086_/Q sky130_fd_sc_hd__dfrtp_4
X_21298_ _15645_/A _21307_/B VGND VGND VPWR VPWR _21304_/B sky130_fd_sc_hd__or2_4
XFILLER_104_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23037_ _23037_/A _22968_/B _22853_/X VGND VGND VPWR VPWR _23037_/X sky130_fd_sc_hd__and3_4
X_20249_ _11865_/X VGND VGND VPWR VPWR _20249_/X sky130_fd_sc_hd__buf_2
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16626__B1 _16368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14810_ _25054_/Q _14810_/B _25055_/Q VGND VGND VPWR VPWR _14811_/B sky130_fd_sc_hd__or3_4
X_15790_ _15758_/A VGND VGND VPWR VPWR _15790_/X sky130_fd_sc_hd__buf_2
X_24988_ _24989_/CLK _24988_/D HRESETn VGND VGND VPWR VPWR _24988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12112__B1 _11834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14741_ _14734_/A _14715_/X _14740_/X VGND VGND VPWR VPWR _14742_/A sky130_fd_sc_hd__a21o_4
X_11953_ _11951_/Y _11944_/X _11952_/X _11944_/X VGND VGND VPWR VPWR _25511_/D sky130_fd_sc_hd__a2bb2o_4
X_23939_ _25154_/CLK _23939_/D HRESETn VGND VGND VPWR VPWR _23939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19550__B _16464_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17460_ _18937_/B VGND VGND VPWR VPWR _18333_/B sky130_fd_sc_hd__inv_2
X_14672_ _19028_/B _19054_/C _19054_/D _19346_/A VGND VGND VPWR VPWR _14672_/X sky130_fd_sc_hd__and4_4
X_11884_ _11884_/A VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__inv_2
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16411_ _15098_/Y _16409_/X _16410_/X _16409_/X VGND VGND VPWR VPWR _24606_/D sky130_fd_sc_hd__a2bb2o_4
X_13623_ _17950_/A _19142_/B _17950_/A _19142_/B VGND VGND VPWR VPWR _14801_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_199_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17391_ _17391_/A _17391_/B VGND VGND VPWR VPWR _17392_/C sky130_fd_sc_hd__nand2_4
XANTENNA__21304__C _21308_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_231_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _25204_/CLK sky130_fd_sc_hd__clkbuf_1
X_19130_ _19130_/A VGND VGND VPWR VPWR _19130_/Y sky130_fd_sc_hd__inv_2
X_16342_ _16341_/Y _16339_/X _16245_/X _16339_/X VGND VGND VPWR VPWR _24630_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13554_ _13552_/Y _25093_/Q _13553_/Y _25099_/Q VGND VGND VPWR VPWR _13563_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12505_ _12263_/Y _12479_/B _12421_/A _12503_/B VGND VGND VPWR VPWR _12505_/X sky130_fd_sc_hd__a211o_4
X_19061_ _19061_/A VGND VGND VPWR VPWR _19061_/X sky130_fd_sc_hd__buf_2
X_16273_ _16273_/A VGND VGND VPWR VPWR _16273_/Y sky130_fd_sc_hd__inv_2
X_13485_ _13484_/X VGND VGND VPWR VPWR _13486_/A sky130_fd_sc_hd__inv_2
XANTENNA__12179__B1 SCLK_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18012_ _18231_/A _18012_/B VGND VGND VPWR VPWR _18012_/X sky130_fd_sc_hd__or2_4
X_15224_ _15075_/C _15221_/X VGND VGND VPWR VPWR _15224_/X sky130_fd_sc_hd__or2_4
X_12436_ _12403_/A _12432_/Y _12436_/C VGND VGND VPWR VPWR _12437_/A sky130_fd_sc_hd__or3_4
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15155_ _15153_/Y _16445_/A _25009_/Q _15154_/Y VGND VGND VPWR VPWR _15155_/X sky130_fd_sc_hd__a2bb2o_4
X_12367_ _12367_/A VGND VGND VPWR VPWR _12997_/C sky130_fd_sc_hd__inv_2
X_14106_ _25229_/Q VGND VGND VPWR VPWR _14128_/C sky130_fd_sc_hd__inv_2
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16865__B1 _16729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12298_ _12424_/A _12261_/Y _12298_/C _12297_/X VGND VGND VPWR VPWR _12299_/B sky130_fd_sc_hd__or4_4
X_15086_ _24591_/Q VGND VGND VPWR VPWR _15086_/Y sky130_fd_sc_hd__inv_2
X_19963_ _21211_/B _19958_/X _19900_/X _19958_/A VGND VGND VPWR VPWR _19963_/X sky130_fd_sc_hd__a2bb2o_4
X_14037_ _14013_/A _14013_/B _14058_/A VGND VGND VPWR VPWR _14037_/Y sky130_fd_sc_hd__o21ai_4
X_18914_ _18914_/A _13757_/A _13754_/X VGND VGND VPWR VPWR _18914_/X sky130_fd_sc_hd__or3_4
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19894_ _23591_/Q VGND VGND VPWR VPWR _19894_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16430__A _16430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18845_ _18841_/X _18842_/X _18843_/X _18844_/X VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__or4_4
XFILLER_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18776_ _18776_/A _18774_/X _18775_/X VGND VGND VPWR VPWR _24146_/D sky130_fd_sc_hd__and3_4
X_15988_ _12219_/Y _15986_/X _15629_/X _15986_/X VGND VGND VPWR VPWR _15988_/X sky130_fd_sc_hd__a2bb2o_4
X_17727_ _17727_/A VGND VGND VPWR VPWR _21675_/A sky130_fd_sc_hd__buf_2
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14939_ _14939_/A VGND VGND VPWR VPWR _14939_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13851__B1 _13806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_41_0_HCLK clkbuf_5_20_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17658_ _17575_/A _17658_/B VGND VGND VPWR VPWR _17658_/X sky130_fd_sc_hd__or2_4
XFILLER_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16609_ HWDATA[9] VGND VGND VPWR VPWR _16609_/X sky130_fd_sc_hd__buf_2
XFILLER_90_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17589_ _17589_/A _17589_/B _17589_/C VGND VGND VPWR VPWR _17589_/X sky130_fd_sc_hd__or3_4
XFILLER_149_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19328_ _23787_/Q VGND VGND VPWR VPWR _19328_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11740__C _11740_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21141__A2 _14229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21511__A _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19259_ _19258_/Y VGND VGND VPWR VPWR _19259_/X sky130_fd_sc_hd__buf_2
X_22270_ _18300_/B _19885_/Y VGND VGND VPWR VPWR _22272_/B sky130_fd_sc_hd__or2_4
XFILLER_157_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21221_ _21280_/A _21220_/Y _24231_/Q _21280_/A VGND VGND VPWR VPWR _21221_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24746__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21152_ _13798_/B _24196_/Q _25175_/Q _12068_/X VGND VGND VPWR VPWR _21153_/B sky130_fd_sc_hd__o22a_4
X_20103_ _20099_/Y _20101_/X _20102_/X _20101_/X VGND VGND VPWR VPWR _20103_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21083_ _21083_/A _21034_/X VGND VGND VPWR VPWR _21083_/X sky130_fd_sc_hd__or2_4
X_20034_ _19900_/A VGND VGND VPWR VPWR _20034_/X sky130_fd_sc_hd__buf_2
X_24911_ _24022_/CLK _24911_/D HRESETn VGND VGND VPWR VPWR _24911_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_247_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24842_ _25425_/CLK _15824_/X HRESETn VGND VGND VPWR VPWR _24842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24773_ _24777_/CLK _24773_/D HRESETn VGND VGND VPWR VPWR _24773_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _24235_/Q _13824_/X VGND VGND VPWR VPWR _21985_/X sky130_fd_sc_hd__or2_4
XFILLER_214_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _23716_/CLK _23724_/D VGND VGND VPWR VPWR _23724_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _24070_/Q VGND VGND VPWR VPWR _20936_/Y sky130_fd_sc_hd__inv_2
XFILLER_242_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _16711_/Y _20854_/X _20863_/X _20866_/X VGND VGND VPWR VPWR _20867_/X sky130_fd_sc_hd__o22a_4
X_23655_ _23654_/CLK _23655_/D VGND VGND VPWR VPWR _19710_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_214_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15595__B1 _11787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22606_ _22563_/X _22605_/X _22145_/C _24871_/Q _22565_/X VGND VGND VPWR VPWR _22606_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20798_ _20797_/Y _20794_/Y _13144_/X VGND VGND VPWR VPWR _20798_/X sky130_fd_sc_hd__o21a_4
X_23586_ _23560_/CLK _19911_/X VGND VGND VPWR VPWR _19909_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17336__A1 _17262_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25325_ _25181_/CLK _25325_/D HRESETn VGND VGND VPWR VPWR _25325_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_210_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22537_ _22506_/X _22510_/X _22516_/Y _22536_/X VGND VGND VPWR VPWR HRDATA[9] sky130_fd_sc_hd__a211o_4
XFILLER_183_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_61_0_HCLK clkbuf_8_61_0_HCLK/A VGND VGND VPWR VPWR _24372_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_155_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13270_ _13417_/A _13270_/B VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__or2_4
X_25256_ _25204_/CLK _13877_/X HRESETn VGND VGND VPWR VPWR _20681_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22468_ _21974_/A VGND VGND VPWR VPWR _22468_/X sky130_fd_sc_hd__buf_2
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12221_ _12210_/X _12214_/X _12221_/C _12221_/D VGND VGND VPWR VPWR _12236_/C sky130_fd_sc_hd__or4_4
X_24207_ _24206_/CLK _24207_/D HRESETn VGND VGND VPWR VPWR _18366_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21419_ _14700_/X _21417_/X _21418_/X VGND VGND VPWR VPWR _21419_/X sky130_fd_sc_hd__and3_4
X_22399_ _21525_/Y _22370_/X _19550_/C _22398_/X VGND VGND VPWR VPWR _22399_/Y sky130_fd_sc_hd__a22oi_4
X_25187_ _25177_/CLK _25187_/D HRESETn VGND VGND VPWR VPWR _13531_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__18836__B2 _18737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24961__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _20981_/A VGND VGND VPWR VPWR _12152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16847__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24138_ _24138_/CLK _18812_/X HRESETn VGND VGND VPWR VPWR _24138_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A VGND VGND VPWR VPWR _12083_/X sky130_fd_sc_hd__buf_2
X_16960_ _16955_/X _16956_/X _16958_/X _16959_/X VGND VGND VPWR VPWR _16961_/D sky130_fd_sc_hd__or4_4
X_24069_ _24503_/CLK _20935_/X HRESETn VGND VGND VPWR VPWR _13659_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_104_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21891__A1_N _12828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22396__A1 _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15911_ _12755_/Y _15908_/X _15632_/X _15908_/X VGND VGND VPWR VPWR _15911_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16891_ _16888_/Y _16889_/X _16890_/X _16889_/X VGND VGND VPWR VPWR _24413_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _24138_/Q VGND VGND VPWR VPWR _18630_/Y sky130_fd_sc_hd__inv_2
X_15842_ _15806_/Y VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__buf_2
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18561_ _18474_/Y _18559_/A VGND VGND VPWR VPWR _18561_/X sky130_fd_sc_hd__or2_4
XFILLER_76_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15773_ _12572_/Y _15772_/X _15636_/X _15772_/X VGND VGND VPWR VPWR _15773_/X sky130_fd_sc_hd__a2bb2o_4
X_12985_ _12853_/Y _12988_/B VGND VGND VPWR VPWR _12985_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13833__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17512_ _17512_/A VGND VGND VPWR VPWR _17569_/B sky130_fd_sc_hd__inv_2
XFILLER_217_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14724_ _21277_/A VGND VGND VPWR VPWR _22237_/A sky130_fd_sc_hd__buf_2
XFILLER_217_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_28_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11936_ _11932_/Y _11935_/X RsRx_S1 _11935_/X VGND VGND VPWR VPWR _25515_/D sky130_fd_sc_hd__a2bb2o_4
X_18492_ _18492_/A _18492_/B _18491_/Y VGND VGND VPWR VPWR _24194_/D sky130_fd_sc_hd__and3_4
XFILLER_33_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17443_ _24332_/Q VGND VGND VPWR VPWR _17443_/Y sky130_fd_sc_hd__inv_2
X_14655_ _18097_/A VGND VGND VPWR VPWR _14656_/A sky130_fd_sc_hd__buf_2
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11867_ _15486_/A VGND VGND VPWR VPWR _11867_/X sky130_fd_sc_hd__buf_2
XFILLER_221_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ _19595_/A _14442_/A VGND VGND VPWR VPWR _13606_/X sky130_fd_sc_hd__or2_4
XFILLER_232_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17374_ _17358_/C _17380_/A VGND VGND VPWR VPWR _17378_/B sky130_fd_sc_hd__or2_4
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14586_ _14593_/A _14582_/Y _14586_/C _14595_/A VGND VGND VPWR VPWR _14586_/X sky130_fd_sc_hd__and4_4
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17327__A1 _17263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11798_ _11796_/Y _11794_/X _11797_/X _11794_/X VGND VGND VPWR VPWR _25543_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22427__A _21604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19113_ _21626_/B _19112_/X _16894_/X _19112_/X VGND VGND VPWR VPWR _23863_/D sky130_fd_sc_hd__a2bb2o_4
X_16325_ _16325_/A VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__buf_2
XANTENNA__21331__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13537_ _13523_/A _13535_/Y _13536_/X _13532_/X VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__a211o_4
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12953__A _12855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16425__A _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22146__B _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19044_ _19037_/A VGND VGND VPWR VPWR _19044_/X sky130_fd_sc_hd__buf_2
XFILLER_146_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16256_ _24661_/Q VGND VGND VPWR VPWR _16256_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13468_ _13468_/A _23613_/Q VGND VGND VPWR VPWR _13469_/C sky130_fd_sc_hd__or2_4
XFILLER_139_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15207_ _15068_/X _15205_/X _15206_/X VGND VGND VPWR VPWR _25038_/D sky130_fd_sc_hd__and3_4
X_12419_ _12403_/A VGND VGND VPWR VPWR _12421_/A sky130_fd_sc_hd__buf_2
X_16187_ _14772_/A _16186_/Y _14769_/X _16186_/Y VGND VGND VPWR VPWR _24685_/D sky130_fd_sc_hd__a2bb2o_4
X_13399_ _13241_/X _13395_/X _13398_/X VGND VGND VPWR VPWR _13399_/X sky130_fd_sc_hd__or3_4
XFILLER_160_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _15137_/Y _16432_/A _15137_/Y _16432_/A VGND VGND VPWR VPWR _15141_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21831__B1 _21697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22162__A _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15069_ _15206_/A _15203_/A VGND VGND VPWR VPWR _15069_/X sky130_fd_sc_hd__or2_4
X_19946_ _19958_/A VGND VGND VPWR VPWR _19946_/X sky130_fd_sc_hd__buf_2
XFILLER_141_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19877_ _21410_/B _19874_/X _19810_/X _19874_/X VGND VGND VPWR VPWR _23598_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18828_ _18621_/X _18828_/B VGND VGND VPWR VPWR _18828_/X sky130_fd_sc_hd__or2_4
XFILLER_95_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18759_ _18759_/A VGND VGND VPWR VPWR _18759_/Y sky130_fd_sc_hd__inv_2
XFILLER_243_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18087__A _18234_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21770_ _21625_/A _21770_/B VGND VGND VPWR VPWR _21770_/X sky130_fd_sc_hd__or2_4
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21225__B _21225_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20721_ _24021_/Q _13137_/B _20725_/B VGND VGND VPWR VPWR _20721_/Y sky130_fd_sc_hd__a21boi_4
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20652_ _17411_/X VGND VGND VPWR VPWR _20669_/C sky130_fd_sc_hd__buf_2
X_23440_ _23441_/CLK _23440_/D VGND VGND VPWR VPWR _23440_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23371_ VGND VGND VPWR VPWR _23371_/HI sda_o_S5 sky130_fd_sc_hd__conb_1
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20583_ _20583_/A VGND VGND VPWR VPWR _23955_/D sky130_fd_sc_hd__inv_2
X_25110_ _23970_/CLK _14536_/X HRESETn VGND VGND VPWR VPWR _25110_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_48_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_97_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22322_ _22321_/X VGND VGND VPWR VPWR _22322_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_19_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22253_ _22027_/A _22253_/B VGND VGND VPWR VPWR _22253_/X sky130_fd_sc_hd__or2_4
X_25041_ _25043_/CLK _15192_/Y HRESETn VGND VGND VPWR VPWR _15002_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24580__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19646__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21204_ _21204_/A _21204_/B _21204_/C VGND VGND VPWR VPWR _21204_/X sky130_fd_sc_hd__and3_4
XANTENNA__20625__A1 _14877_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16829__B1 HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23948__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22184_ _17378_/A _21321_/A _25444_/Q _21081_/A VGND VGND VPWR VPWR _22184_/X sky130_fd_sc_hd__a2bb2o_4
X_21135_ _21135_/A _21135_/B _13781_/A _11718_/B VGND VGND VPWR VPWR _21348_/B sky130_fd_sc_hd__or4_4
XFILLER_132_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15501__B1 HWRITE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16070__A _14423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21066_ _21066_/A _21065_/X VGND VGND VPWR VPWR _21066_/X sky130_fd_sc_hd__or2_4
XFILLER_59_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22800__A _22535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20017_ _20016_/Y VGND VGND VPWR VPWR _20017_/X sky130_fd_sc_hd__buf_2
XFILLER_247_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24825_ _24825_/CLK _24825_/D HRESETn VGND VGND VPWR VPWR _24825_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21889__B1 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12770_ _21035_/A VGND VGND VPWR VPWR _12770_/Y sky130_fd_sc_hd__inv_2
X_24756_ _24756_/CLK _24756_/D HRESETn VGND VGND VPWR VPWR _21715_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21135__B _21135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _21968_/A VGND VGND VPWR VPWR _21968_/X sky130_fd_sc_hd__buf_2
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A VGND VGND VPWR VPWR _11721_/Y sky130_fd_sc_hd__inv_2
X_23707_ _23690_/CLK _23707_/D VGND VGND VPWR VPWR _19554_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20918_/X VGND VGND VPWR VPWR _20924_/B sky130_fd_sc_hd__inv_2
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _24689_/CLK _24687_/D HRESETn VGND VGND VPWR VPWR _21444_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _22093_/A _21899_/B VGND VGND VPWR VPWR _21899_/X sky130_fd_sc_hd__or2_4
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14439_/Y _14435_/X _14409_/X _14428_/A VGND VGND VPWR VPWR _25143_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _23631_/CLK _19759_/X VGND VGND VPWR VPWR _13433_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13869__A _24008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24668__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _25164_/Q _14360_/X _25163_/Q _14365_/X VGND VGND VPWR VPWR _14371_/X sky130_fd_sc_hd__o22a_4
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23569_ _23513_/CLK _23569_/D VGND VGND VPWR VPWR _19953_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12773__A _12773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16245__A _16245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _24712_/Q VGND VGND VPWR VPWR _16110_/Y sky130_fd_sc_hd__inv_2
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13322_/A _13322_/B _13322_/C VGND VGND VPWR VPWR _13323_/C sky130_fd_sc_hd__and3_4
X_25308_ _25494_/CLK _25308_/D HRESETn VGND VGND VPWR VPWR _25308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17090_ _17037_/Y _17088_/X _17089_/Y VGND VGND VPWR VPWR _24403_/D sky130_fd_sc_hd__o21a_4
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16041_ _16040_/Y _16036_/X _15972_/X _16036_/X VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__a2bb2o_4
X_13253_ _13241_/X _13247_/X _13252_/X VGND VGND VPWR VPWR _13253_/X sky130_fd_sc_hd__or3_4
X_25239_ _25246_/CLK _14091_/X HRESETn VGND VGND VPWR VPWR _13999_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_183_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15740__B1 _11783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18460__A _18710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ _12293_/A _12202_/Y _12191_/A _12203_/Y VGND VGND VPWR VPWR _12204_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13184_ _13176_/X _13181_/X _13183_/X VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__o21a_4
X_19800_ _19800_/A VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__buf_2
XFILLER_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12135_ _24115_/Q _12135_/B VGND VGND VPWR VPWR _12136_/B sky130_fd_sc_hd__and2_4
XANTENNA__17076__A _17393_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17992_ _18006_/A VGND VGND VPWR VPWR _18209_/A sky130_fd_sc_hd__buf_2
XFILLER_78_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16943_ _16118_/Y _17751_/A _16118_/Y _17751_/A VGND VGND VPWR VPWR _16943_/X sky130_fd_sc_hd__a2bb2o_4
X_19731_ _19730_/Y _19725_/X _19612_/X _19725_/X VGND VGND VPWR VPWR _23648_/D sky130_fd_sc_hd__a2bb2o_4
X_12066_ _11731_/B VGND VGND VPWR VPWR _19594_/B sky130_fd_sc_hd__inv_2
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23030__A2 _21890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17804__A _17753_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16874_ _20108_/A VGND VGND VPWR VPWR _16874_/X sky130_fd_sc_hd__buf_2
X_19662_ _13329_/B VGND VGND VPWR VPWR _19662_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18993__B1 _18991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15825_ _15758_/A VGND VGND VPWR VPWR _15825_/X sky130_fd_sc_hd__buf_2
X_18613_ _16590_/Y _24147_/Q _16590_/Y _24147_/Q VGND VGND VPWR VPWR _18613_/X sky130_fd_sc_hd__a2bb2o_4
X_19593_ _23692_/Q VGND VGND VPWR VPWR _19593_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20222__A2_N _20219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15756_ HWDATA[13] VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__buf_2
X_18544_ _18540_/B _18550_/B VGND VGND VPWR VPWR _18548_/B sky130_fd_sc_hd__or2_4
XFILLER_206_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12968_ _12952_/C _12952_/D VGND VGND VPWR VPWR _12969_/B sky130_fd_sc_hd__or2_4
XFILLER_80_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14707_ _14695_/Y _14728_/A _14707_/C _14707_/D VGND VGND VPWR VPWR _14707_/X sky130_fd_sc_hd__or4_4
X_11919_ _17711_/B _11889_/A _11911_/X _11918_/Y VGND VGND VPWR VPWR _11919_/X sky130_fd_sc_hd__a211o_4
X_18475_ _18475_/A VGND VGND VPWR VPWR _18484_/B sky130_fd_sc_hd__inv_2
X_15687_ _15920_/B VGND VGND VPWR VPWR _15693_/A sky130_fd_sc_hd__buf_2
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12899_ _12899_/A _12899_/B VGND VGND VPWR VPWR _12901_/B sky130_fd_sc_hd__or2_4
X_17426_ _17426_/A VGND VGND VPWR VPWR _17426_/X sky130_fd_sc_hd__buf_2
X_14638_ _14634_/Y _14637_/Y _14633_/X _14637_/A VGND VGND VPWR VPWR _25087_/D sky130_fd_sc_hd__o22a_4
XFILLER_178_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23260__B _15681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22157__A _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21061__A _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17357_ _17357_/A _17356_/X VGND VGND VPWR VPWR _17380_/A sky130_fd_sc_hd__or2_4
X_14569_ _13561_/Y _14569_/B VGND VGND VPWR VPWR _14570_/B sky130_fd_sc_hd__or2_4
XANTENNA__12683__A _12618_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ _16308_/A VGND VGND VPWR VPWR _16308_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17288_ _17296_/A VGND VGND VPWR VPWR _17288_/X sky130_fd_sc_hd__buf_2
X_19027_ _13628_/A _19142_/B _14668_/A VGND VGND VPWR VPWR _19028_/C sky130_fd_sc_hd__or3_4
X_16239_ _16237_/Y _16235_/X _16238_/X _16235_/X VGND VGND VPWR VPWR _24667_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19466__A _19460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15731__B1 _11766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21798__A1_N _22549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19929_ _19928_/Y _19926_/X _19793_/X _19926_/X VGND VGND VPWR VPWR _19929_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21721__A1_N _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22940_ _22940_/A VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__buf_2
XFILLER_205_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18984__B1 _17430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22871_ _22871_/A _23322_/B VGND VGND VPWR VPWR _22871_/X sky130_fd_sc_hd__or2_4
XFILLER_228_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24610_ _24613_/CLK _16401_/X HRESETn VGND VGND VPWR VPWR _24610_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11762__A _25553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21822_ _21688_/A _21822_/B VGND VGND VPWR VPWR _21822_/X sky130_fd_sc_hd__or2_4
XFILLER_221_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24541_ _24537_/CLK _24541_/D HRESETn VGND VGND VPWR VPWR _16578_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_224_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21753_ _16625_/Y _21588_/X _21591_/A _21752_/X VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__o22a_4
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21886__A3 _22662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20704_ _20724_/A VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__buf_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24472_ _24437_/CLK _24472_/D HRESETn VGND VGND VPWR VPWR _24472_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23088__A2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21684_ _21493_/A _21682_/X _21684_/C VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__and3_4
XANTENNA__14222__B1 _13524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _23400_/CLK _20355_/X VGND VGND VPWR VPWR _23423_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24761__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20635_ _20635_/A VGND VGND VPWR VPWR _20635_/Y sky130_fd_sc_hd__inv_2
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22835__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16065__A _16065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20566_ _20566_/A _18878_/X VGND VGND VPWR VPWR _20566_/Y sky130_fd_sc_hd__nand2_4
X_23354_ _13795_/Y _23354_/B VGND VGND VPWR VPWR _23354_/Y sky130_fd_sc_hd__nor2_4
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22305_ _22430_/A _22305_/B VGND VGND VPWR VPWR _22305_/X sky130_fd_sc_hd__and2_4
XANTENNA__14525__A1 _20609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20497_ _20504_/A _20497_/B _20511_/C VGND VGND VPWR VPWR _20497_/X sky130_fd_sc_hd__and3_4
X_23285_ _23280_/Y _23284_/Y _22868_/X VGND VGND VPWR VPWR _23285_/X sky130_fd_sc_hd__o21a_4
X_25024_ _25018_/CLK _15264_/X HRESETn VGND VGND VPWR VPWR _25024_/Q sky130_fd_sc_hd__dfrtp_4
X_22236_ _22221_/A _22236_/B _22235_/X VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__or3_4
XFILLER_106_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_135_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23654_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_246_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_198_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24674_/CLK sky130_fd_sc_hd__clkbuf_1
X_22167_ _22053_/X _22137_/X _22150_/X _22167_/D VGND VGND VPWR VPWR HRDATA[5] sky130_fd_sc_hd__or4_4
XFILLER_132_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23048__D _23047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21118_ _21082_/X _21083_/X _21100_/X _21112_/X _21117_/X VGND VGND VPWR VPWR _21292_/C
+ sky130_fd_sc_hd__a32o_4
X_22098_ _22228_/A _22093_/X _22094_/X _22095_/X _22097_/X VGND VGND VPWR VPWR _22098_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_87_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13940_ _13940_/A VGND VGND VPWR VPWR _13940_/Y sky130_fd_sc_hd__inv_2
X_21049_ _16280_/A _21105_/B VGND VGND VPWR VPWR _21049_/X sky130_fd_sc_hd__and2_4
XFILLER_75_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23345__B _23313_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13871_ _13871_/A VGND VGND VPWR VPWR _13871_/Y sky130_fd_sc_hd__inv_2
X_15610_ _15608_/Y _15609_/X _11809_/X _15609_/X VGND VGND VPWR VPWR _15610_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16683__A1_N _16682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23242__A1_N _17243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12822_ _12822_/A VGND VGND VPWR VPWR _12912_/A sky130_fd_sc_hd__buf_2
X_24808_ _24812_/CLK _24808_/D HRESETn VGND VGND VPWR VPWR _22875_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16590_ _24536_/Q VGND VGND VPWR VPWR _16590_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15541_ _15540_/Y _15538_/X HADDR[6] _15538_/X VGND VGND VPWR VPWR _24936_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24849__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12753_ _25404_/Q VGND VGND VPWR VPWR _12869_/A sky130_fd_sc_hd__inv_2
X_24739_ _24738_/CLK _16039_/X HRESETn VGND VGND VPWR VPWR _24739_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11702_/A _24233_/Q _13691_/A _11703_/Y VGND VGND VPWR VPWR _11704_/X sky130_fd_sc_hd__o22a_4
X_18260_ _11686_/Y _18258_/X _17433_/X _18258_/X VGND VGND VPWR VPWR _24236_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15472_/A VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__buf_2
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12618_/C _12683_/X VGND VGND VPWR VPWR _12685_/D sky130_fd_sc_hd__or2_4
XANTENNA__14213__B1 _13846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17181_/X _17211_/B _17211_/C _17210_/X VGND VGND VPWR VPWR _17240_/A sky130_fd_sc_hd__or4_4
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14423_/A VGND VGND VPWR VPWR _14423_/X sky130_fd_sc_hd__buf_2
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18191_ _18191_/A _18191_/B _18191_/C VGND VGND VPWR VPWR _18191_/X sky130_fd_sc_hd__and3_4
XANTENNA__22287__B1 _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15961__B1 _15960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _17142_/A _17142_/B VGND VGND VPWR VPWR _17142_/X sky130_fd_sc_hd__or2_4
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ _14347_/Y _14354_/B VGND VGND VPWR VPWR _14359_/B sky130_fd_sc_hd__or2_4
XFILLER_155_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20837__B2 _20836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15310__C _15082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _13207_/X _13304_/X _25336_/Q _13267_/X VGND VGND VPWR VPWR _25336_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_31_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17073_ _17095_/A _17073_/B _17073_/C VGND VGND VPWR VPWR _24407_/D sky130_fd_sc_hd__and3_4
XFILLER_156_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14285_ _21157_/A _14280_/X _13819_/X _14268_/A VGND VGND VPWR VPWR _25190_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22424__B _22424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_94_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16024_ _16019_/A VGND VGND VPWR VPWR _16024_/X sky130_fd_sc_hd__buf_2
X_13236_ _13320_/A VGND VGND VPWR VPWR _13282_/A sky130_fd_sc_hd__buf_2
XFILLER_108_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11847__A _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _13195_/A _23796_/Q VGND VGND VPWR VPWR _13169_/B sky130_fd_sc_hd__or2_4
XFILLER_170_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12118_ _25480_/Q VGND VGND VPWR VPWR _12118_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13098_ _13002_/C _13096_/X _13097_/Y VGND VGND VPWR VPWR _13098_/X sky130_fd_sc_hd__o21a_4
X_17975_ _13613_/A VGND VGND VPWR VPWR _17975_/X sky130_fd_sc_hd__buf_2
XFILLER_111_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22440__A _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_HCLK clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19714_ _19713_/Y _19711_/X _19692_/X _19711_/X VGND VGND VPWR VPWR _23654_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12049_ _25495_/Q VGND VGND VPWR VPWR _12049_/Y sky130_fd_sc_hd__inv_2
X_16926_ _24715_/Q _17787_/A _16102_/Y _16925_/Y VGND VGND VPWR VPWR _16926_/X sky130_fd_sc_hd__o22a_4
X_19645_ _19645_/A VGND VGND VPWR VPWR _21506_/B sky130_fd_sc_hd__inv_2
XANTENNA__20161__A2_N _20156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16857_ _16857_/A VGND VGND VPWR VPWR _16857_/X sky130_fd_sc_hd__buf_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15808_ _15818_/A VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__buf_2
X_16788_ _15037_/Y _16787_/X _16534_/X _16787_/X VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__a2bb2o_4
X_19576_ _22360_/B _19575_/X _11939_/X _19575_/X VGND VGND VPWR VPWR _23700_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22514__A1 _16608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14452__B1 _14427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15739_ _15737_/X _15722_/X _15738_/X _24883_/Q _15720_/X VGND VGND VPWR VPWR _24883_/D
+ sky130_fd_sc_hd__a32o_4
X_18527_ _18527_/A VGND VGND VPWR VPWR _24185_/D sky130_fd_sc_hd__inv_2
XFILLER_206_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14893__A pwm_S6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18458_ _18430_/X _18457_/X VGND VGND VPWR VPWR _18733_/C sky130_fd_sc_hd__or2_4
XFILLER_179_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17409_ _17409_/A VGND VGND VPWR VPWR _17410_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _18388_/Y _18384_/X _24198_/Q _18384_/X VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22817__A2 _22673_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20420_ _20419_/X VGND VGND VPWR VPWR _20420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20351_ _20346_/X VGND VGND VPWR VPWR _20352_/A sky130_fd_sc_hd__inv_2
XANTENNA__23227__C1 _23226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16613__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23070_ _15588_/Y _23140_/B VGND VGND VPWR VPWR _23070_/X sky130_fd_sc_hd__and2_4
XFILLER_161_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20282_ _22207_/B _20279_/X _16870_/X _20279_/X VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__a2bb2o_4
X_22021_ _21936_/A VGND VGND VPWR VPWR _22034_/A sky130_fd_sc_hd__buf_2
XANTENNA__25378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_208_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24532_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22450__B1 _21456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23972_ _24012_/CLK _23972_/D HRESETn VGND VGND VPWR VPWR _14389_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_111_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18957__B1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22923_ _22436_/X _22912_/X _22923_/C _22922_/X VGND VGND VPWR VPWR _22923_/X sky130_fd_sc_hd__or4_4
XFILLER_110_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22854_ _24468_/Q _22854_/B _22853_/X VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__and3_4
XFILLER_232_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21805_ _21493_/A _21803_/X _21804_/X VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__and3_4
XANTENNA__24942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22785_ _22488_/X _22783_/X _21434_/X _24876_/Q _22784_/X VGND VGND VPWR VPWR _22786_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ _24528_/CLK _16624_/X HRESETn VGND VGND VPWR VPWR _16622_/A sky130_fd_sc_hd__dfrtp_4
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21736_ _21736_/A VGND VGND VPWR VPWR _21739_/C sky130_fd_sc_hd__inv_2
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24455_ _24430_/CLK _24455_/D HRESETn VGND VGND VPWR VPWR _15036_/A sky130_fd_sc_hd__dfrtp_4
X_21667_ _21493_/A _21665_/X _21666_/X VGND VGND VPWR VPWR _21667_/X sky130_fd_sc_hd__and3_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23406_ _23582_/CLK _20399_/X VGND VGND VPWR VPWR _23406_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14424__A1_N _14137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13212__A _13212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20618_ _20462_/X _20477_/C _20549_/B VGND VGND VPWR VPWR _20618_/X sky130_fd_sc_hd__o21a_4
X_24386_ _24386_/CLK _17152_/X HRESETn VGND VGND VPWR VPWR _24386_/Q sky130_fd_sc_hd__dfrtp_4
X_21598_ _22768_/A VGND VGND VPWR VPWR _21604_/A sky130_fd_sc_hd__buf_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23337_ _22476_/A _23335_/Y _22479_/A _23336_/Y VGND VGND VPWR VPWR _23338_/B sky130_fd_sc_hd__o22a_4
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20549_ _14543_/A _20549_/B _14024_/X VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__and3_4
XANTENNA__12509__B1 _12403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14070_ _14058_/A _14066_/X _14069_/X VGND VGND VPWR VPWR _25247_/D sky130_fd_sc_hd__o21ai_4
X_23268_ _12790_/Y _21890_/X _16925_/Y _22839_/X VGND VGND VPWR VPWR _23268_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13021_ _13021_/A _13026_/C _13021_/C _13021_/D VGND VGND VPWR VPWR _13022_/A sky130_fd_sc_hd__or4_4
X_25007_ _25002_/CLK _25007_/D HRESETn VGND VGND VPWR VPWR _25007_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22219_ _22227_/A _22219_/B VGND VGND VPWR VPWR _22220_/C sky130_fd_sc_hd__or2_4
XANTENNA__22441__B1 _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23199_ _23199_/A _23119_/B VGND VGND VPWR VPWR _23199_/X sky130_fd_sc_hd__or2_4
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14972_ _14972_/A _14966_/X _14972_/C _14972_/D VGND VGND VPWR VPWR _14993_/B sky130_fd_sc_hd__or4_4
X_17760_ _17861_/A _16916_/Y _17760_/C _17759_/X VGND VGND VPWR VPWR _17761_/D sky130_fd_sc_hd__or4_4
XFILLER_248_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18948__B1 _16791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ _13923_/A _13936_/D _13937_/B _13900_/X VGND VGND VPWR VPWR _13924_/D sky130_fd_sc_hd__or4_4
X_16711_ _24491_/Q VGND VGND VPWR VPWR _16711_/Y sky130_fd_sc_hd__inv_2
X_17691_ _17691_/A VGND VGND VPWR VPWR _17702_/C sky130_fd_sc_hd__buf_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _24518_/Q _16641_/Y _16636_/X VGND VGND VPWR VPWR _16642_/X sky130_fd_sc_hd__o21a_4
X_19430_ _19428_/Y _19429_/X _19383_/X _19429_/X VGND VGND VPWR VPWR _23751_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13854_ _13574_/Y _13852_/X _13812_/X _13852_/X VGND VGND VPWR VPWR _25262_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12805_ _22139_/A VGND VGND VPWR VPWR _12805_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24683__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _16571_/Y _16567_/X _16402_/X _16572_/X VGND VGND VPWR VPWR _24544_/D sky130_fd_sc_hd__a2bb2o_4
X_19361_ _19359_/Y _19360_/X _19226_/X _19360_/X VGND VGND VPWR VPWR _19361_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21604__A _21604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13785_ _19550_/C VGND VGND VPWR VPWR _13804_/C sky130_fd_sc_hd__buf_2
XANTENNA__20507__B1 _20499_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15524_ _15524_/A VGND VGND VPWR VPWR _15524_/Y sky130_fd_sc_hd__inv_2
X_18312_ _21485_/A _18310_/X _18311_/Y VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__o21a_4
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24612__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12736_ _12735_/X VGND VGND VPWR VPWR _25410_/D sky130_fd_sc_hd__inv_2
X_19292_ _23799_/Q VGND VGND VPWR VPWR _21625_/B sky130_fd_sc_hd__inv_2
XFILLER_187_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18243_ _18243_/A VGND VGND VPWR VPWR _18243_/X sky130_fd_sc_hd__buf_2
XFILLER_188_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15455_ _15440_/X VGND VGND VPWR VPWR _15455_/X sky130_fd_sc_hd__buf_2
X_12667_ _12660_/B VGND VGND VPWR VPWR _12671_/B sky130_fd_sc_hd__inv_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _25153_/Q VGND VGND VPWR VPWR _14406_/Y sky130_fd_sc_hd__inv_2
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ _18072_/X _19385_/A VGND VGND VPWR VPWR _18174_/X sky130_fd_sc_hd__or2_4
X_15386_ _15385_/X VGND VGND VPWR VPWR _15386_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12598_ _12589_/X _12598_/B _12594_/X _12597_/X VGND VGND VPWR VPWR _12608_/C sky130_fd_sc_hd__or4_4
XFILLER_184_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22435__A _22401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17125_ _17042_/D _17101_/B _17076_/X _17122_/Y VGND VGND VPWR VPWR _17126_/A sky130_fd_sc_hd__a211o_4
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ _25174_/Q _12172_/X _14336_/Y VGND VGND VPWR VPWR _14337_/X sky130_fd_sc_hd__o21a_4
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17056_ _17086_/D _17086_/B VGND VGND VPWR VPWR _17057_/D sky130_fd_sc_hd__or2_4
XFILLER_116_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14268_ _14268_/A VGND VGND VPWR VPWR _14268_/X sky130_fd_sc_hd__buf_2
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12274__A1_N _12273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23224__A2 _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16007_ _15999_/Y _16006_/X _11752_/X _16006_/X VGND VGND VPWR VPWR _16007_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17439__B1 _16796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23134__A1_N _17305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13219_ _13228_/A VGND VGND VPWR VPWR _13420_/A sky130_fd_sc_hd__buf_2
X_14199_ _14199_/A _14199_/B VGND VGND VPWR VPWR _14204_/A sky130_fd_sc_hd__or2_4
XFILLER_97_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_181_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _25137_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17264__A _17257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_38_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _25066_/CLK sky130_fd_sc_hd__clkbuf_1
X_17958_ _17943_/A _17958_/B VGND VGND VPWR VPWR _17958_/X sky130_fd_sc_hd__or2_4
XFILLER_238_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16909_ _16909_/A VGND VGND VPWR VPWR _17824_/A sky130_fd_sc_hd__inv_2
X_17889_ _17758_/Y _17888_/X _16964_/X VGND VGND VPWR VPWR _17889_/Y sky130_fd_sc_hd__a21oi_4
X_19628_ _23683_/Q VGND VGND VPWR VPWR _19628_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19559_ _23705_/Q VGND VGND VPWR VPWR _19559_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22570_ _22494_/X _22568_/X _21303_/A _24835_/Q _22569_/X VGND VGND VPWR VPWR _22570_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21171__B1 _16192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21521_ _13792_/A VGND VGND VPWR VPWR _22062_/A sky130_fd_sc_hd__buf_2
XFILLER_178_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24240_ _24240_/CLK _18255_/X HRESETn VGND VGND VPWR VPWR _22525_/A sky130_fd_sc_hd__dfrtp_4
X_21452_ _21316_/X VGND VGND VPWR VPWR _22531_/B sky130_fd_sc_hd__buf_2
XFILLER_166_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20403_ _21181_/B _20398_/X _19900_/A _20385_/Y VGND VGND VPWR VPWR _23404_/D sky130_fd_sc_hd__a2bb2o_4
X_21383_ _21383_/A VGND VGND VPWR VPWR _21383_/Y sky130_fd_sc_hd__inv_2
X_24171_ _24171_/CLK _18581_/X HRESETn VGND VGND VPWR VPWR _18414_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12871__A _12609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23122_ _23118_/X _23122_/B VGND VGND VPWR VPWR _23132_/C sky130_fd_sc_hd__and2_4
X_20334_ _21819_/B _20329_/X _20003_/X _20329_/X VGND VGND VPWR VPWR _23431_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16350__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20265_ _13313_/B VGND VGND VPWR VPWR _20265_/Y sky130_fd_sc_hd__inv_2
X_23053_ _23053_/A VGND VGND VPWR VPWR _23119_/B sky130_fd_sc_hd__buf_2
XFILLER_89_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22004_ _22003_/A _21991_/B VGND VGND VPWR VPWR _22004_/X sky130_fd_sc_hd__or2_4
X_20196_ _22219_/B _20193_/X _20105_/X _20193_/X VGND VGND VPWR VPWR _23483_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20985__B1 _14550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20068__A2_N _20065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23955_ _23954_/CLK _23955_/D HRESETn VGND VGND VPWR VPWR _20579_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14948__D _14947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_9_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22906_ _22950_/A _22906_/B _22906_/C VGND VGND VPWR VPWR _22907_/D sky130_fd_sc_hd__and3_4
XFILLER_56_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23886_ _23459_/CLK _19049_/X VGND VGND VPWR VPWR _18189_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22837_ _21293_/X VGND VGND VPWR VPWR _22837_/X sky130_fd_sc_hd__buf_2
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13570_ _25265_/Q _14610_/A _25271_/Q _14581_/A VGND VGND VPWR VPWR _13573_/C sky130_fd_sc_hd__a2bb2o_4
X_25556_ _24732_/CLK _25556_/D HRESETn VGND VGND VPWR VPWR _25556_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22768_ _22768_/A _22768_/B VGND VGND VPWR VPWR _22768_/Y sky130_fd_sc_hd__nor2_4
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A VGND VGND VPWR VPWR _12521_/Y sky130_fd_sc_hd__inv_2
X_24507_ _24073_/CLK _16674_/X HRESETn VGND VGND VPWR VPWR _16671_/A sky130_fd_sc_hd__dfrtp_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21719_ _24620_/Q _21719_/B VGND VGND VPWR VPWR _21719_/X sky130_fd_sc_hd__or2_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15916__B1 _15486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25487_ _25488_/CLK _25487_/D HRESETn VGND VGND VPWR VPWR _12092_/A sky130_fd_sc_hd__dfrtp_4
X_22699_ _22676_/X _22681_/Y _22698_/X VGND VGND VPWR VPWR HRDATA[13] sky130_fd_sc_hd__a21o_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15053_/X _15218_/X VGND VGND VPWR VPWR _15240_/X sky130_fd_sc_hd__or2_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12197_/X _12449_/D VGND VGND VPWR VPWR _12453_/B sky130_fd_sc_hd__or2_4
X_24438_ _24437_/CLK _16829_/X HRESETn VGND VGND VPWR VPWR _14936_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19548__B _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15171_ _15171_/A _15171_/B _15161_/X _15170_/X VGND VGND VPWR VPWR _15171_/X sky130_fd_sc_hd__or4_4
XFILLER_138_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17349__A _17257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12383_ _25370_/Q VGND VGND VPWR VPWR _13011_/A sky130_fd_sc_hd__inv_2
X_24369_ _24372_/CLK _24369_/D HRESETn VGND VGND VPWR VPWR _17310_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14122_ _23968_/Q _14108_/B _25219_/Q VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__or3_4
XFILLER_126_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25143__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14053_ _14028_/A _14027_/D _14053_/C _14027_/B VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__or4_4
X_18930_ _18928_/Y _18929_/X _16894_/X _18929_/X VGND VGND VPWR VPWR _23927_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13004_ _12351_/Y _13004_/B _13115_/A _13088_/A VGND VGND VPWR VPWR _13004_/X sky130_fd_sc_hd__or4_4
X_18861_ _18861_/A _18861_/B _18861_/C _18860_/X VGND VGND VPWR VPWR _18861_/X sky130_fd_sc_hd__or4_4
XFILLER_67_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_254_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _24003_/CLK sky130_fd_sc_hd__clkbuf_1
X_17812_ _17751_/A _17815_/B VGND VGND VPWR VPWR _17813_/C sky130_fd_sc_hd__or2_4
XFILLER_239_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17084__A _17393_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18792_ _18685_/Y _18791_/X VGND VGND VPWR VPWR _18809_/B sky130_fd_sc_hd__or2_4
XANTENNA__14501__A _25119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15998__A3 _15933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14955_ _25014_/Q _14953_/Y _15282_/A _14954_/Y VGND VGND VPWR VPWR _14960_/B sky130_fd_sc_hd__a2bb2o_4
X_17743_ _17743_/A _17743_/B _17736_/X _17742_/X VGND VGND VPWR VPWR _17743_/X sky130_fd_sc_hd__or4_4
XANTENNA__24864__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18908__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _13936_/D VGND VGND VPWR VPWR _13927_/B sky130_fd_sc_hd__buf_2
XFILLER_235_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17812__A _17751_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14886_ _14873_/B _14880_/X _14881_/Y VGND VGND VPWR VPWR _14886_/Y sky130_fd_sc_hd__a21oi_4
X_17674_ _17588_/A _17693_/A VGND VGND VPWR VPWR _17674_/X sky130_fd_sc_hd__or2_4
XANTENNA__14407__B1 _14248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19413_ _14665_/Y _19143_/B _19346_/C VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__or3_4
X_13837_ _13553_/Y _13834_/X _11827_/X _13834_/X VGND VGND VPWR VPWR _13837_/X sky130_fd_sc_hd__a2bb2o_4
X_16625_ _16625_/A VGND VGND VPWR VPWR _16625_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12956__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11860__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _24550_/Q VGND VGND VPWR VPWR _16556_/Y sky130_fd_sc_hd__inv_2
X_19344_ _19343_/Y _19338_/X _19254_/X _19324_/Y VGND VGND VPWR VPWR _23781_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13768_ _13768_/A VGND VGND VPWR VPWR _13768_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12719_ _12623_/C _12722_/B _12662_/X VGND VGND VPWR VPWR _12719_/Y sky130_fd_sc_hd__a21oi_4
X_15507_ _11736_/A VGND VGND VPWR VPWR _15507_/Y sky130_fd_sc_hd__inv_2
X_16487_ _24576_/Q VGND VGND VPWR VPWR _16487_/Y sky130_fd_sc_hd__inv_2
X_19275_ _19275_/A VGND VGND VPWR VPWR _21243_/B sky130_fd_sc_hd__inv_2
XANTENNA__15907__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13699_ _11688_/Y _13699_/B VGND VGND VPWR VPWR _13700_/B sky130_fd_sc_hd__or2_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15438_ _13959_/X _15438_/B _15438_/C _14255_/B VGND VGND VPWR VPWR _15444_/A sky130_fd_sc_hd__or4_4
X_18226_ _18063_/A _18226_/B _18226_/C VGND VGND VPWR VPWR _18227_/C sky130_fd_sc_hd__and3_4
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16580__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19649__B2 _19624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24345__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15369_ _15139_/Y _15360_/X VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__or2_4
X_18157_ _18090_/A _18157_/B VGND VGND VPWR VPWR _18157_/X sky130_fd_sc_hd__or2_4
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17108_ _17108_/A VGND VGND VPWR VPWR _17108_/Y sky130_fd_sc_hd__inv_2
X_18088_ _17954_/A _18079_/X _18088_/C VGND VGND VPWR VPWR _18088_/X sky130_fd_sc_hd__and3_4
XFILLER_171_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17039_ _24394_/Q VGND VGND VPWR VPWR _17042_/B sky130_fd_sc_hd__inv_2
X_20050_ _20050_/A VGND VGND VPWR VPWR _20050_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16635__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23740_ _23794_/CLK _23740_/D VGND VGND VPWR VPWR _17965_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_227_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15536__A2_N _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _20952_/A VGND VGND VPWR VPWR _20952_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16399__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23669_/CLK _23671_/D VGND VGND VPWR VPWR _13397_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20883_/A VGND VGND VPWR VPWR _20883_/X sky130_fd_sc_hd__buf_2
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16338__A _16338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25410_ _25410_/CLK _25410_/D HRESETn VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23133__B2 _22924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11770__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22622_ _12851_/A _22678_/B _22621_/X VGND VGND VPWR VPWR _22622_/X sky130_fd_sc_hd__o21a_4
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25341_ _25368_/CLK _25341_/D HRESETn VGND VGND VPWR VPWR _13003_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22553_ _24057_/Q _21320_/A _13139_/A _21322_/X VGND VGND VPWR VPWR _22553_/Y sky130_fd_sc_hd__a22oi_4
X_21504_ _21473_/A VGND VGND VPWR VPWR _21668_/A sky130_fd_sc_hd__buf_2
XFILLER_194_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25272_ _25103_/CLK _25272_/D HRESETn VGND VGND VPWR VPWR _25272_/Q sky130_fd_sc_hd__dfrtp_4
X_22484_ _22157_/C VGND VGND VPWR VPWR _22484_/X sky130_fd_sc_hd__buf_2
XFILLER_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _24295_/CLK _24223_/D HRESETn VGND VGND VPWR VPWR _17733_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_148_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21447__A1 _15565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21435_ _11744_/X VGND VGND VPWR VPWR _22578_/B sky130_fd_sc_hd__buf_2
XANTENNA__21447__B2 _22530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16073__A _14427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18312__A1 _21485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24154_ _23976_/CLK _18745_/X HRESETn VGND VGND VPWR VPWR _24154_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21366_ _12109_/A _17448_/B _21362_/X _21577_/A _21365_/X VGND VGND VPWR VPWR _21366_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__16323__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22803__A _16689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23105_ _12216_/Y _22444_/X _22730_/X _12330_/Y _22858_/X VGND VGND VPWR VPWR _23105_/X
+ sky130_fd_sc_hd__o32a_4
X_20317_ _23437_/Q VGND VGND VPWR VPWR _21469_/B sky130_fd_sc_hd__inv_2
XFILLER_190_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24085_ _24966_/CLK _20544_/X HRESETn VGND VGND VPWR VPWR _24085_/Q sky130_fd_sc_hd__dfrtp_4
X_21297_ _21877_/B VGND VGND VPWR VPWR _21307_/B sky130_fd_sc_hd__buf_2
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23036_ _15158_/A _22849_/X VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__or2_4
XFILLER_89_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20248_ _20234_/Y VGND VGND VPWR VPWR _20248_/X sky130_fd_sc_hd__buf_2
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20179_ _23489_/Q VGND VGND VPWR VPWR _20179_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_21_0_HCLK clkbuf_7_10_0_HCLK/X VGND VGND VPWR VPWR _24272_/CLK sky130_fd_sc_hd__clkbuf_1
X_24987_ _24989_/CLK _24987_/D HRESETn VGND VGND VPWR VPWR _24987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_84_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _25368_/CLK sky130_fd_sc_hd__clkbuf_1
X_14740_ _14735_/X _14739_/Y _14732_/Y VGND VGND VPWR VPWR _14740_/X sky130_fd_sc_hd__a21o_4
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ _19636_/A VGND VGND VPWR VPWR _11952_/X sky130_fd_sc_hd__buf_2
X_23938_ _24012_/CLK _23938_/D HRESETn VGND VGND VPWR VPWR _23938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19550__C _19550_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14671_ _25079_/Q VGND VGND VPWR VPWR _19346_/A sky130_fd_sc_hd__buf_2
X_11883_ _25524_/Q _11897_/A _11884_/A VGND VGND VPWR VPWR _11883_/Y sky130_fd_sc_hd__a21oi_4
X_23869_ _23871_/CLK _19096_/X VGND VGND VPWR VPWR _13442_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_199_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16248__A _16248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12776__A _25381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ HWDATA[21] VGND VGND VPWR VPWR _16410_/X sky130_fd_sc_hd__buf_2
X_13622_ _25076_/Q VGND VGND VPWR VPWR _19142_/B sky130_fd_sc_hd__buf_2
X_17390_ _17363_/A _17390_/B _17389_/Y VGND VGND VPWR VPWR _24348_/D sky130_fd_sc_hd__and3_4
XFILLER_199_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ _24630_/Q VGND VGND VPWR VPWR _16341_/Y sky130_fd_sc_hd__inv_2
X_13553_ _25271_/Q VGND VGND VPWR VPWR _13553_/Y sky130_fd_sc_hd__inv_2
X_25539_ _25539_/CLK _25539_/D HRESETn VGND VGND VPWR VPWR _11811_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12504_ _12501_/A _12500_/B _12504_/C VGND VGND VPWR VPWR _25443_/D sky130_fd_sc_hd__and3_4
X_19060_ _19060_/A VGND VGND VPWR VPWR _19060_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16272_ _16271_/Y _16269_/X _15483_/X _16269_/X VGND VGND VPWR VPWR _24655_/D sky130_fd_sc_hd__a2bb2o_4
X_13484_ _12109_/C _12080_/X _13484_/C _13484_/D VGND VGND VPWR VPWR _13484_/X sky130_fd_sc_hd__or4_4
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15223_ _14912_/X _15223_/B VGND VGND VPWR VPWR _15223_/X sky130_fd_sc_hd__or2_4
X_18011_ _18098_/A VGND VGND VPWR VPWR _18231_/A sky130_fd_sc_hd__buf_2
XANTENNA__12179__B2 _12168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21438__A1 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12435_ _12297_/X _12400_/B _12261_/Y VGND VGND VPWR VPWR _12436_/C sky130_fd_sc_hd__o21a_4
XANTENNA__22635__B1 _22431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ _24613_/Q VGND VGND VPWR VPWR _15154_/Y sky130_fd_sc_hd__inv_2
X_12366_ _13063_/B _24842_/Q _25361_/Q _12317_/Y VGND VGND VPWR VPWR _12369_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20110__B2 _20109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14105_ scl_oen_o_S4 _20996_/B _20419_/B VGND VGND VPWR VPWR _14116_/B sky130_fd_sc_hd__and3_4
XFILLER_154_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15085_ _15322_/A _24616_/Q _15322_/A _24616_/Q VGND VGND VPWR VPWR _15085_/X sky130_fd_sc_hd__a2bb2o_4
X_19962_ _19962_/A VGND VGND VPWR VPWR _21211_/B sky130_fd_sc_hd__inv_2
X_12297_ _12292_/X _12296_/X VGND VGND VPWR VPWR _12297_/X sky130_fd_sc_hd__or2_4
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14036_ _14003_/Y _14030_/X _14556_/B VGND VGND VPWR VPWR _14060_/A sky130_fd_sc_hd__a21o_4
X_18913_ _14706_/A VGND VGND VPWR VPWR _20149_/B sky130_fd_sc_hd__buf_2
XFILLER_106_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19893_ _21806_/B _19888_/X _19639_/X _19888_/X VGND VGND VPWR VPWR _23592_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17814__B1 _16952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15327__A _15324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11855__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18844_ _24554_/Q _24133_/Q _16544_/Y _18689_/B VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__o22a_4
XFILLER_228_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12580__A2_N _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18775_ _18694_/Y _18773_/A VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__or2_4
X_15987_ _12213_/Y _15983_/X _15767_/X _15986_/X VGND VGND VPWR VPWR _24761_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ _21936_/A VGND VGND VPWR VPWR _17727_/A sky130_fd_sc_hd__buf_2
XFILLER_236_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14938_ _15188_/A VGND VGND VPWR VPWR _15182_/A sky130_fd_sc_hd__inv_2
XANTENNA__21064__A _21032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17657_ _17644_/X VGND VGND VPWR VPWR _17658_/B sky130_fd_sc_hd__inv_2
XFILLER_223_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14869_ _14854_/X _14868_/Y _24961_/Q _14820_/X VGND VGND VPWR VPWR _25051_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19319__B1 _19184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16608_ _24529_/Q VGND VGND VPWR VPWR _16608_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17588_ _17588_/A _17588_/B _17537_/Y _17587_/Y VGND VGND VPWR VPWR _17589_/C sky130_fd_sc_hd__or4_4
XFILLER_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19327_ _19322_/Y _19325_/X _19326_/X _19325_/X VGND VGND VPWR VPWR _19327_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16539_ _24556_/Q VGND VGND VPWR VPWR _16539_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11740__D _11740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19258_ _19258_/A VGND VGND VPWR VPWR _19258_/Y sky130_fd_sc_hd__inv_2
X_18209_ _18209_/A _18209_/B VGND VGND VPWR VPWR _18211_/B sky130_fd_sc_hd__or2_4
X_19189_ _19346_/A _19143_/B _19028_/C VGND VGND VPWR VPWR _19189_/X sky130_fd_sc_hd__or3_4
XFILLER_191_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11917__A1 _11890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _21220_/A VGND VGND VPWR VPWR _21220_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21151_ _13526_/Y _21031_/X _21577_/B _21150_/Y VGND VGND VPWR VPWR _21155_/A sky130_fd_sc_hd__a211o_4
XFILLER_171_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20102_ _20102_/A VGND VGND VPWR VPWR _20102_/X sky130_fd_sc_hd__buf_2
X_21082_ _21082_/A VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__buf_2
XANTENNA__24786__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20033_ _20033_/A VGND VGND VPWR VPWR _20033_/Y sky130_fd_sc_hd__inv_2
X_24910_ _24020_/CLK _15617_/X HRESETn VGND VGND VPWR VPWR _15616_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14779__C _13599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24715__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17281__A1 _17270_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24841_ _24889_/CLK _15827_/X HRESETn VGND VGND VPWR VPWR _24841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_1_0_HCLK_A clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19558__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17452__A _19139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24772_ _24792_/CLK _24772_/D HRESETn VGND VGND VPWR VPWR _22910_/A sky130_fd_sc_hd__dfrtp_4
X_21984_ _19550_/C _21983_/X VGND VGND VPWR VPWR _21984_/Y sky130_fd_sc_hd__nand2_4
XFILLER_215_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ _23716_/CLK _23723_/D VGND VGND VPWR VPWR _23723_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _20927_/X _20934_/Y _24506_/Q _20931_/X VGND VGND VPWR VPWR _20935_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16068__A _24727_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23654_/CLK _23654_/D VGND VGND VPWR VPWR _19713_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20864_/Y _20859_/Y _20865_/X VGND VGND VPWR VPWR _20866_/X sky130_fd_sc_hd__o21a_4
XFILLER_241_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22605_ _22605_/A _21104_/B VGND VGND VPWR VPWR _22605_/X sky130_fd_sc_hd__or2_4
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23560_/CLK _23585_/D VGND VGND VPWR VPWR _23585_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ _20797_/A VGND VGND VPWR VPWR _20797_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25324_ _25181_/CLK _25324_/D HRESETn VGND VGND VPWR VPWR _13497_/A sky130_fd_sc_hd__dfrtp_4
X_22536_ _22536_/A _22536_/B _22529_/Y _22535_/Y VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__or4_4
X_25255_ _25200_/CLK _25255_/D HRESETn VGND VGND VPWR VPWR _25255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22467_ _16284_/X _22467_/B VGND VGND VPWR VPWR _22480_/A sky130_fd_sc_hd__nor2_4
XFILLER_154_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12220_ _12218_/A _22418_/A _12218_/Y _12219_/Y VGND VGND VPWR VPWR _12221_/D sky130_fd_sc_hd__o22a_4
X_24206_ _24206_/CLK _24206_/D HRESETn VGND VGND VPWR VPWR _24206_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13220__A _13420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21418_ _14765_/X _21418_/B VGND VGND VPWR VPWR _21418_/X sky130_fd_sc_hd__or2_4
XANTENNA__18297__B1 _17710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25186_ _25177_/CLK _25186_/D HRESETn VGND VGND VPWR VPWR _14296_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22398_ _22237_/A _22377_/Y _22384_/Y _22391_/Y _22397_/Y VGND VGND VPWR VPWR _22398_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22533__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12151_ _12136_/A _12136_/B _12150_/Y VGND VGND VPWR VPWR _20981_/A sky130_fd_sc_hd__o21a_4
X_24137_ _24160_/CLK _24137_/D HRESETn VGND VGND VPWR VPWR _24137_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21840__A1 _21833_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21349_ _21348_/X VGND VGND VPWR VPWR _21731_/A sky130_fd_sc_hd__buf_2
XANTENNA__23348__B _23345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12082_ _12081_/X VGND VGND VPWR VPWR _12083_/A sky130_fd_sc_hd__inv_2
X_24068_ _24503_/CLK _20932_/X HRESETn VGND VGND VPWR VPWR _13659_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15910_ _12784_/Y _15908_/X _15629_/X _15908_/X VGND VGND VPWR VPWR _15910_/X sky130_fd_sc_hd__a2bb2o_4
X_23019_ _22950_/A _23014_/X _23018_/X VGND VGND VPWR VPWR _23020_/D sky130_fd_sc_hd__and3_4
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16890_ _19803_/A VGND VGND VPWR VPWR _16890_/X sky130_fd_sc_hd__buf_2
XANTENNA__20988__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15841_ _12305_/Y _15838_/X _15632_/X _15838_/X VGND VGND VPWR VPWR _24831_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17362__A _17362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18560_ _18474_/A _18560_/B VGND VGND VPWR VPWR _18562_/B sky130_fd_sc_hd__or2_4
XFILLER_206_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23083__B _23080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ _12984_/A _12984_/B _12983_/Y VGND VGND VPWR VPWR _25375_/D sky130_fd_sc_hd__and3_4
X_15772_ _15772_/A VGND VGND VPWR VPWR _15772_/X sky130_fd_sc_hd__buf_2
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20159__B2 _20156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14699__A2_N _14761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17511_ _17511_/A VGND VGND VPWR VPWR _17579_/A sky130_fd_sc_hd__inv_2
X_11935_ _11934_/X VGND VGND VPWR VPWR _11935_/X sky130_fd_sc_hd__buf_2
X_14723_ _14723_/A VGND VGND VPWR VPWR _21277_/A sky130_fd_sc_hd__buf_2
XFILLER_245_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18491_ _18490_/A _18490_/B VGND VGND VPWR VPWR _18491_/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14654_ _13613_/A VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__inv_2
X_17442_ _21567_/A _17441_/X _16861_/X _17441_/X VGND VGND VPWR VPWR _24333_/D sky130_fd_sc_hd__a2bb2o_4
X_11866_ _11865_/X VGND VGND VPWR VPWR _15486_/A sky130_fd_sc_hd__buf_2
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16783__B1 _16609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ _21031_/A _13821_/B _13822_/A _13786_/A VGND VGND VPWR VPWR _14442_/A sky130_fd_sc_hd__or4_4
XFILLER_221_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21612__A _21263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585_ _14563_/Y _14566_/X _14583_/X _25103_/Q _14584_/Y VGND VGND VPWR VPWR _14585_/X
+ sky130_fd_sc_hd__a32o_4
X_17373_ _17372_/X VGND VGND VPWR VPWR _17373_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21659__B2 _22549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ HWDATA[18] VGND VGND VPWR VPWR _11797_/X sky130_fd_sc_hd__buf_2
XPHY_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19112_ _19099_/Y VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__buf_2
XANTENNA__25244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13536_ _13536_/A _25306_/Q VGND VGND VPWR VPWR _13536_/X sky130_fd_sc_hd__and2_4
X_16324_ _24636_/Q VGND VGND VPWR VPWR _16324_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16535__B1 _16534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16255_ _16254_/Y _16251_/X _15905_/X _16251_/X VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__a2bb2o_4
X_19043_ _18157_/B VGND VGND VPWR VPWR _19043_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13467_ _13371_/A _13467_/B VGND VGND VPWR VPWR _13467_/X sky130_fd_sc_hd__or2_4
X_15206_ _15206_/A _15203_/X VGND VGND VPWR VPWR _15206_/X sky130_fd_sc_hd__or2_4
X_12418_ _12398_/A _12418_/B _12417_/X VGND VGND VPWR VPWR _25465_/D sky130_fd_sc_hd__and3_4
XFILLER_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16186_ _16185_/X VGND VGND VPWR VPWR _16186_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23281__B1 _12555_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13398_ _13290_/X _13398_/B _13397_/X VGND VGND VPWR VPWR _13398_/X sky130_fd_sc_hd__and3_4
XANTENNA__22443__A _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15137_ _24993_/Q VGND VGND VPWR VPWR _15137_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12349_ _12310_/X _12349_/B _12349_/C _12348_/X VGND VGND VPWR VPWR _12391_/A sky130_fd_sc_hd__or4_4
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14849__B1 _25202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22162__B _22155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15068_ _15293_/A VGND VGND VPWR VPWR _15068_/X sky130_fd_sc_hd__buf_2
X_19945_ _18290_/X VGND VGND VPWR VPWR _19958_/A sky130_fd_sc_hd__inv_2
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14019_ _14058_/A _14008_/X _14062_/C VGND VGND VPWR VPWR _14553_/A sky130_fd_sc_hd__or3_4
XFILLER_96_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19876_ _19876_/A VGND VGND VPWR VPWR _21410_/B sky130_fd_sc_hd__inv_2
X_18827_ _18749_/A _18824_/B _18826_/Y VGND VGND VPWR VPWR _24132_/D sky130_fd_sc_hd__and3_4
XFILLER_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18758_ _18696_/D _18753_/B _18740_/X _18755_/B VGND VGND VPWR VPWR _18759_/A sky130_fd_sc_hd__a211o_4
XFILLER_67_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17709_ _17708_/X VGND VGND VPWR VPWR _17709_/Y sky130_fd_sc_hd__inv_2
X_18689_ _18689_/A _18689_/B _18689_/C VGND VGND VPWR VPWR _18690_/D sky130_fd_sc_hd__or3_4
XFILLER_24_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20720_ _20720_/A VGND VGND VPWR VPWR _20720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16774__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21522__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20651_ _17402_/A _17402_/B VGND VGND VPWR VPWR _20651_/Y sky130_fd_sc_hd__nand2_4
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15520__A _15503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23370_ VGND VGND VPWR VPWR _23370_/HI sda_o_S4 sky130_fd_sc_hd__conb_1
X_20582_ _14439_/Y _20574_/X _20565_/X _20581_/X VGND VGND VPWR VPWR _20583_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16526__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22321_ _14382_/Y _21861_/A _14483_/Y _21375_/A VGND VGND VPWR VPWR _22321_/X sky130_fd_sc_hd__o22a_4
XFILLER_176_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13040__A _13049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25040_ _25030_/CLK _15197_/X HRESETn VGND VGND VPWR VPWR _15195_/A sky130_fd_sc_hd__dfrtp_4
X_22252_ _22260_/A _22252_/B VGND VGND VPWR VPWR _22252_/X sky130_fd_sc_hd__or2_4
XANTENNA__24967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21203_ _21211_/A _20055_/Y VGND VGND VPWR VPWR _21204_/C sky130_fd_sc_hd__or2_4
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22183_ _22183_/A _22178_/Y _22181_/Y _22182_/X VGND VGND VPWR VPWR _22183_/X sky130_fd_sc_hd__or4_4
XANTENNA__16351__A _24626_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21134_ _17450_/B VGND VGND VPWR VPWR _21134_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21065_ _21064_/X VGND VGND VPWR VPWR _21065_/X sky130_fd_sc_hd__buf_2
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20016_ _20016_/A VGND VGND VPWR VPWR _20016_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23184__A _22897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24824_ _24824_/CLK _15853_/X HRESETn VGND VGND VPWR VPWR _21024_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24755_ _24765_/CLK _24755_/D HRESETn VGND VGND VPWR VPWR _21544_/A sky130_fd_sc_hd__dfrtp_4
X_21967_ _21967_/A VGND VGND VPWR VPWR _21968_/A sky130_fd_sc_hd__buf_2
XFILLER_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _17456_/A VGND VGND VPWR VPWR _14385_/A sky130_fd_sc_hd__buf_2
X_23706_ _23703_/CLK _23706_/D VGND VGND VPWR VPWR _23706_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _13672_/X _13658_/X VGND VGND VPWR VPWR _20918_/X sky130_fd_sc_hd__or2_4
X_24686_ _24726_/CLK _16176_/X HRESETn VGND VGND VPWR VPWR _21069_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16765__B1 _16417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _21263_/A VGND VGND VPWR VPWR _22093_/A sky130_fd_sc_hd__buf_2
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_158_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _24119_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22528__A _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23637_ _23631_/CLK _23637_/D VGND VGND VPWR VPWR _13465_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _20849_/A VGND VGND VPWR VPWR _20849_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _14364_/X _14368_/X _12085_/A _14369_/X VGND VGND VPWR VPWR _14370_/X sky130_fd_sc_hd__o22a_4
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23568_ _23799_/CLK _23568_/D VGND VGND VPWR VPWR _23568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13421_/A _13321_/B VGND VGND VPWR VPWR _13322_/C sky130_fd_sc_hd__or2_4
X_25307_ _25062_/CLK _25307_/D HRESETn VGND VGND VPWR VPWR _13547_/A sky130_fd_sc_hd__dfstp_4
X_22519_ _12032_/Y _13484_/D _12101_/Y _12081_/B VGND VGND VPWR VPWR _22519_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _23516_/CLK _20154_/X VGND VGND VPWR VPWR _20153_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16040_ _24738_/Q VGND VGND VPWR VPWR _16040_/Y sky130_fd_sc_hd__inv_2
X_13252_ _13197_/A _13252_/B _13251_/X VGND VGND VPWR VPWR _13252_/X sky130_fd_sc_hd__and3_4
X_25238_ _25246_/CLK _25238_/D HRESETn VGND VGND VPWR VPWR _25238_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ _23196_/A VGND VGND VPWR VPWR _12203_/Y sky130_fd_sc_hd__inv_2
X_13183_ _13416_/A VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__buf_2
X_25169_ _24121_/CLK _25169_/D HRESETn VGND VGND VPWR VPWR _25169_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24637__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _24113_/Q _12134_/B VGND VGND VPWR VPWR _12135_/B sky130_fd_sc_hd__and2_4
XFILLER_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17991_ _18097_/A VGND VGND VPWR VPWR _17991_/X sky130_fd_sc_hd__buf_2
XFILLER_145_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13503__B1 _13481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19730_ _13368_/B VGND VGND VPWR VPWR _19730_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _11734_/B VGND VGND VPWR VPWR _13542_/C sky130_fd_sc_hd__buf_2
X_16942_ _16143_/Y _17762_/A _16143_/Y _17762_/A VGND VGND VPWR VPWR _16942_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19661_ _19658_/Y _19653_/X _19659_/X _19660_/X VGND VGND VPWR VPWR _19661_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16873_ _16871_/Y _16868_/X _16872_/X _16868_/X VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18188__A _13639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18612_ _18605_/X _18612_/B _18612_/C _18611_/X VGND VGND VPWR VPWR _18643_/A sky130_fd_sc_hd__or4_4
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15824_ _12350_/Y _15821_/X _11800_/X _15821_/X VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__a2bb2o_4
X_19592_ _21194_/B _19587_/X _19501_/X _19574_/Y VGND VGND VPWR VPWR _19592_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18543_ _18543_/A _18543_/B VGND VGND VPWR VPWR _18550_/B sky130_fd_sc_hd__or2_4
XANTENNA__16851__A1_N _14925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_54_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12967_ _12967_/A VGND VGND VPWR VPWR _25381_/D sky130_fd_sc_hd__inv_2
X_15755_ _15737_/X _15751_/X _15754_/X _24874_/Q _15749_/X VGND VGND VPWR VPWR _15755_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _11918_/A VGND VGND VPWR VPWR _11918_/Y sky130_fd_sc_hd__inv_2
X_14706_ _14706_/A _14695_/B VGND VGND VPWR VPWR _14707_/D sky130_fd_sc_hd__and2_4
X_18474_ _18474_/A VGND VGND VPWR VPWR _18474_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12898_ _12900_/B VGND VGND VPWR VPWR _12899_/B sky130_fd_sc_hd__inv_2
X_15686_ _15701_/A VGND VGND VPWR VPWR _15686_/X sky130_fd_sc_hd__buf_2
XANTENNA__22438__A _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ _17424_/X _14232_/B VGND VGND VPWR VPWR _17426_/A sky130_fd_sc_hd__nor2_4
XANTENNA__21342__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11849_ _25530_/Q VGND VGND VPWR VPWR _11849_/Y sky130_fd_sc_hd__inv_2
X_14637_ _14637_/A VGND VGND VPWR VPWR _14637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12964__A _12855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14568_/A VGND VGND VPWR VPWR _14605_/A sky130_fd_sc_hd__inv_2
X_17356_ _17255_/D _17391_/B VGND VGND VPWR VPWR _17356_/X sky130_fd_sc_hd__or2_4
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16307_ _16304_/Y _16305_/X _16306_/X _16305_/X VGND VGND VPWR VPWR _24643_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13519_ _13518_/Y _13516_/X _11862_/X _13516_/X VGND VGND VPWR VPWR _25315_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14499_ _14499_/A VGND VGND VPWR VPWR _14499_/Y sky130_fd_sc_hd__inv_2
X_17287_ _17242_/X _17285_/X _17287_/C VGND VGND VPWR VPWR _24375_/D sky130_fd_sc_hd__and3_4
XFILLER_146_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19026_ _23892_/Q VGND VGND VPWR VPWR _19026_/Y sky130_fd_sc_hd__inv_2
X_16238_ _16238_/A VGND VGND VPWR VPWR _16238_/X sky130_fd_sc_hd__buf_2
XFILLER_173_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17267__A _17245_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _21709_/A VGND VGND VPWR VPWR _16169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16171__A _21531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18276__A3 _13481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22901__A _22171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19928_ _23579_/Q VGND VGND VPWR VPWR _19928_/Y sky130_fd_sc_hd__inv_2
X_19859_ _25285_/Q VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__buf_2
XFILLER_217_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18098__A _18098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22870_ _22832_/X _22836_/X _22870_/C _22869_/X VGND VGND VPWR VPWR HRDATA[17] sky130_fd_sc_hd__or4_4
XANTENNA__21236__B _21046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21821_ _21687_/A _19914_/Y VGND VGND VPWR VPWR _21821_/X sky130_fd_sc_hd__or2_4
XFILLER_209_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24540_ _24537_/CLK _24540_/D HRESETn VGND VGND VPWR VPWR _24540_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_221_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13035__A _13049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21752_ _16542_/Y _21752_/B VGND VGND VPWR VPWR _21752_/X sky130_fd_sc_hd__and2_4
XFILLER_169_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16747__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21740__B1 _24588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _20702_/X VGND VGND VPWR VPWR _20703_/Y sky130_fd_sc_hd__inv_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24471_ _24437_/CLK _24471_/D HRESETn VGND VGND VPWR VPWR _24471_/Q sky130_fd_sc_hd__dfrtp_4
X_21683_ _21688_/A _21683_/B VGND VGND VPWR VPWR _21684_/C sky130_fd_sc_hd__or2_4
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14222__B2 _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23422_ _24206_/CLK _23422_/D VGND VGND VPWR VPWR _23422_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20634_ _15479_/Y _20623_/X _20680_/A _20633_/X VGND VGND VPWR VPWR _20635_/A sky130_fd_sc_hd__a211o_4
XFILLER_196_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23353_ _23353_/A VGND VGND VPWR VPWR _23353_/Y sky130_fd_sc_hd__inv_2
X_20565_ _20564_/X VGND VGND VPWR VPWR _20565_/X sky130_fd_sc_hd__buf_2
XFILLER_164_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22304_ _21431_/X _22302_/X _22303_/X _24866_/Q _22558_/A VGND VGND VPWR VPWR _22305_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23284_ _23283_/X VGND VGND VPWR VPWR _23284_/Y sky130_fd_sc_hd__inv_2
X_20496_ _24088_/Q _20520_/A VGND VGND VPWR VPWR _20511_/C sky130_fd_sc_hd__and2_4
XFILLER_152_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22083__A _22390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25023_ _25023_/CLK _25023_/D HRESETn VGND VGND VPWR VPWR _25023_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22599__A2 _22596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22235_ _22235_/A _22235_/B _22234_/X VGND VGND VPWR VPWR _22235_/X sky130_fd_sc_hd__and3_4
XANTENNA__24730__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22166_ _22152_/X _22165_/X VGND VGND VPWR VPWR _22167_/D sky130_fd_sc_hd__and2_4
XANTENNA__18672__B1 _16625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21117_ _17251_/A _21113_/X _21116_/X VGND VGND VPWR VPWR _21117_/X sky130_fd_sc_hd__o21a_4
X_22097_ _22385_/A _19866_/Y _22209_/A VGND VGND VPWR VPWR _22097_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22530__B _22530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21048_ _15673_/A VGND VGND VPWR VPWR _21048_/X sky130_fd_sc_hd__buf_2
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15238__B1 _15208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13870_ _13869_/X VGND VGND VPWR VPWR _13870_/X sky130_fd_sc_hd__buf_2
XFILLER_207_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20782__A1 _22934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12821_ _25388_/Q VGND VGND VPWR VPWR _12822_/A sky130_fd_sc_hd__inv_2
X_24807_ _24856_/CLK _15893_/X HRESETn VGND VGND VPWR VPWR _24807_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12364__A2_N _24848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22999_ _12293_/Y _22998_/X _16909_/A _22924_/X VGND VGND VPWR VPWR _22999_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12752_ _12851_/A _22605_/A _12851_/A _22605_/A VGND VGND VPWR VPWR _12752_/X sky130_fd_sc_hd__a2bb2o_4
X_15540_ _21135_/B VGND VGND VPWR VPWR _15540_/Y sky130_fd_sc_hd__inv_2
X_24738_ _24738_/CLK _16041_/X HRESETn VGND VGND VPWR VPWR _24738_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _24233_/Q VGND VGND VPWR VPWR _11703_/Y sky130_fd_sc_hd__inv_2
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _15471_/A _14232_/B VGND VGND VPWR VPWR _15472_/A sky130_fd_sc_hd__nor2_4
X_12683_ _12618_/D _12674_/X VGND VGND VPWR VPWR _12683_/X sky130_fd_sc_hd__or2_4
X_24669_ _24552_/CLK _24669_/D HRESETn VGND VGND VPWR VPWR _16231_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12784__A _22428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ HWDATA[6] VGND VGND VPWR VPWR _14423_/A sky130_fd_sc_hd__buf_2
X_17210_ _17202_/X _17204_/X _17210_/C _17210_/D VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__or4_4
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12379__A2_N _12377_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18158_/A _23878_/Q VGND VGND VPWR VPWR _18191_/C sky130_fd_sc_hd__or2_4
XANTENNA__13599__B _13599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24889__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12775__A1 _12773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _14352_/X VGND VGND VPWR VPWR _14354_/B sky130_fd_sc_hd__buf_2
X_17141_ _16987_/Y _17157_/A VGND VGND VPWR VPWR _17142_/B sky130_fd_sc_hd__or2_4
XFILLER_7_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24818__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13304_ _13209_/X _13285_/X _13303_/X _25337_/Q _11974_/X VGND VGND VPWR VPWR _13304_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17072_/A _17072_/B VGND VGND VPWR VPWR _17073_/C sky130_fd_sc_hd__or2_4
X_14284_ _14284_/A VGND VGND VPWR VPWR _21157_/A sky130_fd_sc_hd__inv_2
XFILLER_144_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12302__A2_N _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13235_ _13356_/A _18942_/A VGND VGND VPWR VPWR _13238_/B sky130_fd_sc_hd__or2_4
X_16023_ _24745_/Q VGND VGND VPWR VPWR _16023_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _13451_/A VGND VGND VPWR VPWR _13197_/A sky130_fd_sc_hd__buf_2
XFILLER_3_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22721__A _16338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12117_ _12140_/A _12111_/X _11842_/X _12116_/X VGND VGND VPWR VPWR _12117_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13097_ _13002_/C _13096_/X _13040_/X VGND VGND VPWR VPWR _13097_/Y sky130_fd_sc_hd__a21oi_4
X_17974_ _14794_/A VGND VGND VPWR VPWR _18227_/A sky130_fd_sc_hd__buf_2
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19713_ _19713_/A VGND VGND VPWR VPWR _19713_/Y sky130_fd_sc_hd__inv_2
X_12048_ _12047_/Y _12043_/X _25495_/Q _12043_/X VGND VGND VPWR VPWR _12048_/X sky130_fd_sc_hd__a2bb2o_4
X_16925_ _17787_/A VGND VGND VPWR VPWR _16925_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18415__B1 _16259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15229__B1 _15183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19644_ _21695_/B _19642_/X _19643_/X _19642_/X VGND VGND VPWR VPWR _23679_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16856_ _24423_/Q VGND VGND VPWR VPWR _16856_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15807_ _15806_/Y VGND VGND VPWR VPWR _15818_/A sky130_fd_sc_hd__buf_2
X_19575_ _19574_/Y VGND VGND VPWR VPWR _19575_/X sky130_fd_sc_hd__buf_2
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16787_ _16782_/A VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__buf_2
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13999_ _13999_/A _13999_/B _13999_/C _13999_/D VGND VGND VPWR VPWR _14000_/C sky130_fd_sc_hd__or4_4
X_18526_ _18828_/B _18523_/B _18525_/X VGND VGND VPWR VPWR _18527_/A sky130_fd_sc_hd__or3_4
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15738_ HWDATA[23] VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__buf_2
XFILLER_222_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18457_ _18438_/X _18457_/B _18451_/X _18456_/X VGND VGND VPWR VPWR _18457_/X sky130_fd_sc_hd__or4_4
X_15669_ _15652_/Y _15664_/X _15656_/X _20830_/A _15668_/X VGND VGND VPWR VPWR _15669_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_141_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23642_/CLK sky130_fd_sc_hd__clkbuf_1
X_17408_ _23999_/Q _17408_/B VGND VGND VPWR VPWR _17409_/A sky130_fd_sc_hd__or2_4
X_18388_ _24199_/Q VGND VGND VPWR VPWR _18388_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12766__B2 _23162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17339_ _17341_/B VGND VGND VPWR VPWR _17340_/B sky130_fd_sc_hd__inv_2
XANTENNA__24559__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20350_ _23424_/Q VGND VGND VPWR VPWR _20350_/Y sky130_fd_sc_hd__inv_2
X_19009_ _19006_/Y _19004_/X _19008_/X _19004_/X VGND VGND VPWR VPWR _23899_/D sky130_fd_sc_hd__a2bb2o_4
X_20281_ _23451_/Q VGND VGND VPWR VPWR _22207_/B sky130_fd_sc_hd__inv_2
XANTENNA__18249__A3 _16241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22020_ _22265_/A VGND VGND VPWR VPWR _22036_/A sky130_fd_sc_hd__buf_2
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22450__B2 _22449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17725__A _21210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17209__A1 _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17209__B2 _17389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23971_ _25106_/CLK _20616_/X HRESETn VGND VGND VPWR VPWR _23971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11773__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22922_ _22787_/X _22919_/Y _22881_/X _22921_/X VGND VGND VPWR VPWR _22922_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22753__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18957__B2 _18952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22853_ _21589_/B VGND VGND VPWR VPWR _22853_/X sky130_fd_sc_hd__buf_2
XFILLER_71_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21804_ _21497_/A _20312_/Y VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__or2_4
X_22784_ _21436_/X VGND VGND VPWR VPWR _22784_/X sky130_fd_sc_hd__buf_2
XFILLER_25_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21713__B1 _24863_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24523_ _24523_/CLK _16626_/X HRESETn VGND VGND VPWR VPWR _16625_/A sky130_fd_sc_hd__dfrtp_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21735_ _21734_/Y _21161_/X _15482_/Y _21370_/X VGND VGND VPWR VPWR _21736_/A sky130_fd_sc_hd__o22a_4
XFILLER_240_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17610__D _17610_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ _24613_/CLK _16797_/X HRESETn VGND VGND VPWR VPWR _24454_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_240_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21666_ _21468_/X _21666_/B VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__or2_4
XANTENNA__24982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23405_ _23534_/CLK _20401_/X VGND VGND VPWR VPWR _20400_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_196_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20617_ _20465_/X _20473_/B _20549_/B VGND VGND VPWR VPWR _23970_/D sky130_fd_sc_hd__o21a_4
XFILLER_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24385_ _24386_/CLK _17154_/X HRESETn VGND VGND VPWR VPWR _24385_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17145__B1 _17065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24911__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21597_ _21597_/A VGND VGND VPWR VPWR _22768_/A sky130_fd_sc_hd__buf_2
XFILLER_165_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16804__A _16552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22525__B _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23336_/A _16552_/A VGND VGND VPWR VPWR _23336_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20548_ _17429_/A _20548_/B VGND VGND VPWR VPWR _23973_/D sky130_fd_sc_hd__and2_4
XFILLER_4_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12509__A1 _12273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23267_ _23093_/A _23267_/B _23266_/X VGND VGND VPWR VPWR _23267_/X sky130_fd_sc_hd__and3_4
X_20479_ _20437_/A VGND VGND VPWR VPWR _20479_/X sky130_fd_sc_hd__buf_2
XFILLER_180_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13020_ _13020_/A VGND VGND VPWR VPWR _25370_/D sky130_fd_sc_hd__inv_2
X_25006_ _25002_/CLK _25006_/D HRESETn VGND VGND VPWR VPWR _25006_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22218_ _22210_/A _22218_/B VGND VGND VPWR VPWR _22218_/X sky130_fd_sc_hd__or2_4
XFILLER_152_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22441__A1 _16354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23198_ _23117_/A _23197_/X VGND VGND VPWR VPWR _23198_/X sky130_fd_sc_hd__and2_4
XANTENNA__22541__A _22541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22149_ _21714_/A _22140_/X _22145_/X _22148_/X VGND VGND VPWR VPWR _22149_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17635__A _17567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14971_ _15243_/A _24434_/Q _14969_/Y _24434_/Q VGND VGND VPWR VPWR _14972_/D sky130_fd_sc_hd__a2bb2o_4
X_16710_ _16708_/Y _16704_/X _16613_/X _16709_/X VGND VGND VPWR VPWR _16710_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25088__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13922_ _13902_/A VGND VGND VPWR VPWR _13924_/B sky130_fd_sc_hd__inv_2
XFILLER_120_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17690_ _17504_/Y _17674_/X VGND VGND VPWR VPWR _17690_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16959__B1 _16169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16641_ _16640_/X VGND VGND VPWR VPWR _16641_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23372__A _23356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13853_ _13581_/Y _13848_/X _13809_/X _13852_/X VGND VGND VPWR VPWR _13853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17370__A _17364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12804_ _21432_/A VGND VGND VPWR VPWR _12804_/Y sky130_fd_sc_hd__inv_2
X_19360_ _19353_/A VGND VGND VPWR VPWR _19360_/X sky130_fd_sc_hd__buf_2
XANTENNA__23091__B _22954_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16572_ _16584_/A VGND VGND VPWR VPWR _16572_/X sky130_fd_sc_hd__buf_2
X_13784_ _13828_/C VGND VGND VPWR VPWR _19550_/C sky130_fd_sc_hd__buf_2
XFILLER_188_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18311_ _18308_/X VGND VGND VPWR VPWR _18311_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15523_ _15522_/Y _15520_/X HADDR[13] _15520_/X VGND VGND VPWR VPWR _15523_/X sky130_fd_sc_hd__a2bb2o_4
X_12735_ _12590_/Y _12712_/B _12733_/B _12662_/X VGND VGND VPWR VPWR _12735_/X sky130_fd_sc_hd__a211o_4
X_19291_ _21770_/B _19286_/X _16890_/X _19286_/X VGND VGND VPWR VPWR _23800_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18242_ _18241_/Y VGND VGND VPWR VPWR _18243_/A sky130_fd_sc_hd__buf_2
X_12666_ _12636_/A _12666_/B _12665_/Y VGND VGND VPWR VPWR _25430_/D sky130_fd_sc_hd__and3_4
X_15454_ _13951_/B _15446_/X _15441_/X _13951_/A _15453_/X VGND VGND VPWR VPWR _24975_/D
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_214_0_HCLK clkbuf_8_214_0_HCLK/A VGND VGND VPWR VPWR _24425_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _14402_/Y _14403_/X _14404_/X _14393_/X VGND VGND VPWR VPWR _25154_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18832__A1_N _16510_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _17973_/X _18172_/X _24249_/Q _18031_/X VGND VGND VPWR VPWR _24249_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24652__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12588_/A _12595_/Y _12596_/Y _12593_/A VGND VGND VPWR VPWR _12597_/X sky130_fd_sc_hd__a2bb2o_4
X_15385_ _15139_/Y _15360_/X _15324_/X _15383_/B VGND VGND VPWR VPWR _15385_/X sky130_fd_sc_hd__a211o_4
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22435__B _22435_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17106_/A _17120_/B _17123_/X VGND VGND VPWR VPWR _17124_/X sky130_fd_sc_hd__and3_4
XFILLER_156_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ _14335_/X VGND VGND VPWR VPWR _14336_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23209__B1 _16910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14267_ _21726_/B _14232_/B VGND VGND VPWR VPWR _14268_/A sky130_fd_sc_hd__nor2_4
X_17055_ _17132_/A _17129_/A _17055_/C VGND VGND VPWR VPWR _17086_/B sky130_fd_sc_hd__or3_4
XFILLER_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18847__A1_N _24579_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13218_ _13212_/A VGND VGND VPWR VPWR _13228_/A sky130_fd_sc_hd__buf_2
X_16006_ _16005_/X VGND VGND VPWR VPWR _16006_/X sky130_fd_sc_hd__buf_2
X_14198_ _14385_/A _16190_/B _16378_/C _16378_/D VGND VGND VPWR VPWR _14199_/B sky130_fd_sc_hd__or4_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22432__B2 _21322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20361__A1_N _20360_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13149_ _23386_/Q _20696_/B VGND VGND VPWR VPWR _13149_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21067__A _22694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17957_ _17941_/A _17955_/X _17956_/X VGND VGND VPWR VPWR _17957_/X sky130_fd_sc_hd__and3_4
XFILLER_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22196__B1 _21565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ _22574_/A _17861_/C _16110_/Y _24289_/Q VGND VGND VPWR VPWR _16913_/B sky130_fd_sc_hd__a2bb2o_4
X_17888_ _16929_/Y _17891_/B VGND VGND VPWR VPWR _17888_/X sky130_fd_sc_hd__or2_4
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19627_ _19622_/Y _19625_/X _19626_/X _19625_/X VGND VGND VPWR VPWR _23684_/D sky130_fd_sc_hd__a2bb2o_4
X_16839_ _16853_/A VGND VGND VPWR VPWR _16839_/X sky130_fd_sc_hd__buf_2
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15622__B1 _11831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19558_ _19556_/Y _19552_/X _19421_/X _19557_/X VGND VGND VPWR VPWR _23706_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22499__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17711__C _21704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_24_0_HCLK clkbuf_5_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18509_ _24190_/Q _18513_/B VGND VGND VPWR VPWR _18509_/X sky130_fd_sc_hd__or2_4
X_19489_ _19483_/Y VGND VGND VPWR VPWR _19489_/X sky130_fd_sc_hd__buf_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21520_ _21519_/X VGND VGND VPWR VPWR _21520_/X sky130_fd_sc_hd__buf_2
XANTENNA__12855__C _12855_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21710__A3 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22626__A _16432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21530__A _22721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21451_ _21451_/A _21450_/X VGND VGND VPWR VPWR _21451_/X sky130_fd_sc_hd__or2_4
XANTENNA__24393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20402_ _23404_/Q VGND VGND VPWR VPWR _21181_/B sky130_fd_sc_hd__inv_2
X_24170_ _24169_/CLK _24170_/D HRESETn VGND VGND VPWR VPWR _18418_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21382_ _13802_/A _21382_/B _21382_/C VGND VGND VPWR VPWR _21383_/A sky130_fd_sc_hd__or3_4
XANTENNA__15136__A2_N _15134_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23121_ _23052_/X _23119_/X _22986_/X _24885_/Q _23120_/X VGND VGND VPWR VPWR _23122_/B
+ sky130_fd_sc_hd__a32o_4
X_20333_ _23431_/Q VGND VGND VPWR VPWR _21819_/B sky130_fd_sc_hd__inv_2
X_23052_ _21430_/X VGND VGND VPWR VPWR _23052_/X sky130_fd_sc_hd__buf_2
XFILLER_150_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18627__B1 _16612_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20264_ _20262_/Y _20258_/X _19772_/X _20263_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22003_ _22003_/A _21991_/B VGND VGND VPWR VPWR _22003_/X sky130_fd_sc_hd__and2_4
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20195_ _20195_/A VGND VGND VPWR VPWR _22219_/B sky130_fd_sc_hd__inv_2
XANTENNA__20959__A1_N _20836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_106_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23954_ _23954_/CLK _23954_/D HRESETn VGND VGND VPWR VPWR _18881_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22905_ _14922_/A _22541_/A _22542_/A _22904_/X VGND VGND VPWR VPWR _22906_/C sky130_fd_sc_hd__a211o_4
XFILLER_217_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23885_ _23885_/CLK _19051_/X VGND VGND VPWR VPWR _19050_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22836_ _22836_/A _22836_/B _22835_/X VGND VGND VPWR VPWR _22836_/X sky130_fd_sc_hd__and3_4
XFILLER_232_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22767_ _21295_/A _22765_/X _22121_/X _22766_/X VGND VGND VPWR VPWR _22768_/B sky130_fd_sc_hd__o22a_4
X_25555_ _24732_/CLK _11756_/X HRESETn VGND VGND VPWR VPWR _11754_/A sky130_fd_sc_hd__dfrtp_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18563__C1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12520_ _12623_/C _24871_/Q _12623_/C _24871_/Q VGND VGND VPWR VPWR _12520_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21718_ _21126_/B VGND VGND VPWR VPWR _22289_/A sky130_fd_sc_hd__buf_2
X_24506_ _24503_/CLK _24506_/D HRESETn VGND VGND VPWR VPWR _24506_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25486_ _24112_/CLK _12096_/X HRESETn VGND VGND VPWR VPWR _12094_/A sky130_fd_sc_hd__dfrtp_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22698_ _16284_/X _22687_/Y _22689_/Y _22693_/Y _22697_/Y VGND VGND VPWR VPWR _22698_/X
+ sky130_fd_sc_hd__a2111o_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12222_/Y _12449_/X _12450_/Y VGND VGND VPWR VPWR _25457_/D sky130_fd_sc_hd__o21a_4
X_21649_ _21611_/X _21647_/X _21649_/C VGND VGND VPWR VPWR _21649_/X sky130_fd_sc_hd__and3_4
X_24437_ _24437_/CLK _24437_/D HRESETn VGND VGND VPWR VPWR _14922_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16534__A _14423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15170_ _15170_/A _15165_/X _15166_/X _15169_/X VGND VGND VPWR VPWR _15170_/X sky130_fd_sc_hd__or4_4
XANTENNA__24063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12382_ _12381_/Y _24828_/Q _13003_/A _12353_/Y VGND VGND VPWR VPWR _12382_/X sky130_fd_sc_hd__a2bb2o_4
X_24368_ _24639_/CLK _24368_/D HRESETn VGND VGND VPWR VPWR _17231_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_44_0_HCLK clkbuf_7_22_0_HCLK/X VGND VGND VPWR VPWR _23445_/CLK sky130_fd_sc_hd__clkbuf_1
X_14121_ _25228_/Q VGND VGND VPWR VPWR _14121_/Y sky130_fd_sc_hd__inv_2
X_23319_ _24784_/Q _22669_/B VGND VGND VPWR VPWR _23319_/X sky130_fd_sc_hd__or2_4
X_24299_ _25528_/CLK _24299_/D HRESETn VGND VGND VPWR VPWR _24299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14052_ _14052_/A VGND VGND VPWR VPWR _14059_/B sky130_fd_sc_hd__inv_2
XFILLER_180_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22271__A _22271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14989__A _25019_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _13003_/A VGND VGND VPWR VPWR _13115_/A sky130_fd_sc_hd__inv_2
XANTENNA__25269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18860_ _16517_/Y _18693_/A _16517_/Y _18693_/A VGND VGND VPWR VPWR _18860_/X sky130_fd_sc_hd__a2bb2o_4
X_17811_ _17802_/X VGND VGND VPWR VPWR _17815_/B sky130_fd_sc_hd__inv_2
X_18791_ _18690_/D _18791_/B VGND VGND VPWR VPWR _18791_/X sky130_fd_sc_hd__or2_4
XFILLER_153_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17742_ _21509_/A _17741_/X _21509_/A _17741_/X VGND VGND VPWR VPWR _17742_/X sky130_fd_sc_hd__a2bb2o_4
X_14954_ _14954_/A VGND VGND VPWR VPWR _14954_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18397__A2 _17280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13905_ _13923_/A VGND VGND VPWR VPWR _13927_/A sky130_fd_sc_hd__inv_2
XFILLER_208_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17673_ _17588_/B _17672_/X VGND VGND VPWR VPWR _17693_/A sky130_fd_sc_hd__or2_4
X_14885_ _14885_/A VGND VGND VPWR VPWR _14885_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19412_ _19412_/A VGND VGND VPWR VPWR _19412_/Y sky130_fd_sc_hd__inv_2
X_16624_ _16622_/Y _16618_/X _16364_/X _16623_/X VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__a2bb2o_4
X_13836_ _13555_/Y _13834_/X _11822_/X _13834_/X VGND VGND VPWR VPWR _25272_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19343_ _18209_/B VGND VGND VPWR VPWR _19343_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16555_ _16550_/Y _16554_/X _16385_/X _16554_/X VGND VGND VPWR VPWR _24551_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24833__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _25284_/Q _13767_/B VGND VGND VPWR VPWR _13768_/A sky130_fd_sc_hd__and2_4
XANTENNA__14229__A _14229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20113__A2_N _20109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15506_ _16190_/B _15503_/X HADDR[20] _15503_/X VGND VGND VPWR VPWR _15506_/X sky130_fd_sc_hd__a2bb2o_4
X_12718_ _12623_/D _12718_/B VGND VGND VPWR VPWR _12722_/B sky130_fd_sc_hd__or2_4
X_19274_ _21391_/B _19271_/X _16897_/X _19271_/X VGND VGND VPWR VPWR _19274_/X sky130_fd_sc_hd__a2bb2o_4
X_16486_ _16485_/Y _16483_/X _16309_/X _16483_/X VGND VGND VPWR VPWR _16486_/X sky130_fd_sc_hd__a2bb2o_4
X_13698_ _13698_/A _13698_/B VGND VGND VPWR VPWR _13699_/B sky130_fd_sc_hd__or2_4
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18225_ _18129_/A _19024_/A VGND VGND VPWR VPWR _18226_/C sky130_fd_sc_hd__or2_4
X_15437_ _15437_/A _15436_/Y VGND VGND VPWR VPWR _15438_/B sky130_fd_sc_hd__or2_4
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12649_ _12642_/A _12647_/X _12657_/A _12644_/B VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__a211o_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18156_ _13639_/X _18148_/X _18155_/X VGND VGND VPWR VPWR _18156_/X sky130_fd_sc_hd__and3_4
XANTENNA__24083__D _20479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15368_ _15367_/X VGND VGND VPWR VPWR _25001_/D sky130_fd_sc_hd__inv_2
XFILLER_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17107_ _17016_/Y _17101_/X _17076_/X _17104_/B VGND VGND VPWR VPWR _17108_/A sky130_fd_sc_hd__a211o_4
X_14319_ _25182_/Q _14311_/X _25181_/Q _14316_/X VGND VGND VPWR VPWR _14319_/X sky130_fd_sc_hd__o22a_4
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18087_ _18234_/A _18082_/X _18087_/C VGND VGND VPWR VPWR _18088_/C sky130_fd_sc_hd__or3_4
X_15299_ _24483_/Q VGND VGND VPWR VPWR _15299_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17038_ _17037_/Y _17088_/A VGND VGND VPWR VPWR _17057_/C sky130_fd_sc_hd__or2_4
XANTENNA__23277__A _21879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20967__B2 _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18989_ _18988_/Y _18986_/X _18969_/X _18986_/X VGND VGND VPWR VPWR _23905_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15843__B1 _15636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20951_ _20927_/X _20950_/X _16664_/A _20931_/X VGND VGND VPWR VPWR _24073_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23670_ _23669_/CLK _23670_/D VGND VGND VPWR VPWR _13429_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ _20904_/A VGND VGND VPWR VPWR _20883_/A sky130_fd_sc_hd__buf_2
XFILLER_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22621_ _17864_/A _22443_/A _12287_/A _22447_/A VGND VGND VPWR VPWR _22621_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24574__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21144__A1 _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22341__B1 _21565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25340_ _25365_/CLK _13126_/Y HRESETn VGND VGND VPWR VPWR _12320_/A sky130_fd_sc_hd__dfrtp_4
X_22552_ _21321_/X VGND VGND VPWR VPWR _22677_/B sky130_fd_sc_hd__buf_2
XANTENNA__24503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16449__A2_N _16446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16020__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21503_ _21808_/A _21501_/X _21502_/X VGND VGND VPWR VPWR _21503_/X sky130_fd_sc_hd__and3_4
X_25271_ _25103_/CLK _13837_/X HRESETn VGND VGND VPWR VPWR _25271_/Q sky130_fd_sc_hd__dfrtp_4
X_22483_ _22483_/A _23322_/B VGND VGND VPWR VPWR _22483_/X sky130_fd_sc_hd__or2_4
XFILLER_194_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24222_ _24295_/CLK _18295_/X HRESETn VGND VGND VPWR VPWR _24222_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21434_ _22986_/A VGND VGND VPWR VPWR _21434_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_3_0_HCLK clkbuf_7_1_0_HCLK/X VGND VGND VPWR VPWR _23441_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_148_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24153_ _24145_/CLK _18748_/Y HRESETn VGND VGND VPWR VPWR _24153_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21365_ _13504_/B _21363_/X _12108_/B _21364_/X VGND VGND VPWR VPWR _21365_/X sky130_fd_sc_hd__o22a_4
XFILLER_238_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23104_ _22837_/X _23095_/Y _23099_/Y _23103_/X VGND VGND VPWR VPWR _23112_/C sky130_fd_sc_hd__a211o_4
X_20316_ _21666_/B _20315_/X _20007_/X _20315_/X VGND VGND VPWR VPWR _23438_/D sky130_fd_sc_hd__a2bb2o_4
X_24084_ _24966_/CLK _24084_/D HRESETn VGND VGND VPWR VPWR _20540_/B sky130_fd_sc_hd__dfrtp_4
X_21296_ _21322_/A VGND VGND VPWR VPWR _21296_/X sky130_fd_sc_hd__buf_2
XANTENNA__22091__A _22390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23035_ _23035_/A VGND VGND VPWR VPWR _23035_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20247_ _20247_/A VGND VGND VPWR VPWR _20247_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20178_ _20176_/Y _20172_/X _20108_/X _20177_/X VGND VGND VPWR VPWR _23490_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15834__B1 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13218__A _13212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19025__B1 _18999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24986_ _24989_/CLK _24986_/D HRESETn VGND VGND VPWR VPWR _24986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11951_ _19639_/A VGND VGND VPWR VPWR _11951_/Y sky130_fd_sc_hd__inv_2
X_23937_ _24095_/CLK _25118_/Q HRESETn VGND VGND VPWR VPWR _23937_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11961__A _19643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11882_ _17711_/A _11881_/X VGND VGND VPWR VPWR _11884_/A sky130_fd_sc_hd__or2_4
X_14670_ _14670_/A VGND VGND VPWR VPWR _19054_/C sky130_fd_sc_hd__buf_2
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23868_ _23628_/CLK _23868_/D VGND VGND VPWR VPWR _23868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13621_ _18023_/A VGND VGND VPWR VPWR _17950_/A sky130_fd_sc_hd__buf_2
X_22819_ _16733_/A _22819_/B _22818_/X VGND VGND VPWR VPWR _22824_/C sky130_fd_sc_hd__and3_4
XANTENNA__23133__A1_N _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23799_/CLK _23799_/D VGND VGND VPWR VPWR _23799_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16340_ _16338_/Y _16333_/X _16241_/X _16339_/X VGND VGND VPWR VPWR _16340_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _25265_/Q VGND VGND VPWR VPWR _13552_/Y sky130_fd_sc_hd__inv_2
X_25538_ _24732_/CLK _11819_/X HRESETn VGND VGND VPWR VPWR _11816_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12820__B1 _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21170__A _21170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12503_ _12503_/A _12503_/B VGND VGND VPWR VPWR _12504_/C sky130_fd_sc_hd__or2_4
X_13483_ _25329_/Q VGND VGND VPWR VPWR _13483_/Y sky130_fd_sc_hd__inv_2
X_16271_ _24655_/Q VGND VGND VPWR VPWR _16271_/Y sky130_fd_sc_hd__inv_2
X_25469_ _25380_/CLK _25469_/D HRESETn VGND VGND VPWR VPWR _12188_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18010_ _18127_/A _18010_/B _18010_/C VGND VGND VPWR VPWR _18016_/B sky130_fd_sc_hd__and3_4
XFILLER_173_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12434_ _12398_/A _12425_/B _12433_/X VGND VGND VPWR VPWR _25461_/D sky130_fd_sc_hd__and3_4
X_15222_ _15221_/X VGND VGND VPWR VPWR _15223_/B sky130_fd_sc_hd__inv_2
XFILLER_200_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12365_ _25357_/Q VGND VGND VPWR VPWR _13063_/B sky130_fd_sc_hd__inv_2
X_15153_ _15153_/A VGND VGND VPWR VPWR _15153_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22713__B _21855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14104_ _20995_/B VGND VGND VPWR VPWR _20996_/B sky130_fd_sc_hd__inv_2
XFILLER_5_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15084_ _15321_/A VGND VGND VPWR VPWR _15322_/A sky130_fd_sc_hd__inv_2
X_19961_ _19960_/Y _19958_/X _19646_/X _19958_/X VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__a2bb2o_4
X_12296_ _12296_/A _12296_/B _12296_/C _12295_/X VGND VGND VPWR VPWR _12296_/X sky130_fd_sc_hd__or4_4
XFILLER_113_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22399__B1 _19550_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12841__A1_N _25401_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14035_ _14034_/X VGND VGND VPWR VPWR _14556_/B sky130_fd_sc_hd__inv_2
X_18912_ _23932_/Q VGND VGND VPWR VPWR _18912_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19892_ _23592_/Q VGND VGND VPWR VPWR _21806_/B sky130_fd_sc_hd__inv_2
XFILLER_79_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21329__B _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18843_ _24560_/Q _24139_/Q _16527_/Y _18799_/B VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19016__B1 _18969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18774_ _18657_/X _18773_/Y VGND VGND VPWR VPWR _18774_/X sky130_fd_sc_hd__or2_4
X_15986_ _15945_/Y VGND VGND VPWR VPWR _15986_/X sky130_fd_sc_hd__buf_2
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17725_ _21210_/A VGND VGND VPWR VPWR _21936_/A sky130_fd_sc_hd__buf_2
XFILLER_209_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14937_ _25032_/Q _14936_/A _14935_/X _14936_/Y VGND VGND VPWR VPWR _14937_/X sky130_fd_sc_hd__o22a_4
XFILLER_208_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11871__A _14248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17656_ _17641_/A _17649_/X _17656_/C VGND VGND VPWR VPWR _17656_/X sky130_fd_sc_hd__and3_4
XFILLER_236_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14868_ _14868_/A VGND VGND VPWR VPWR _14868_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17261__C _17322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16607_ _16606_/Y _16604_/X _16349_/X _16604_/X VGND VGND VPWR VPWR _24530_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13819_ _16729_/A VGND VGND VPWR VPWR _13819_/X sky130_fd_sc_hd__buf_2
X_17587_ _24296_/Q VGND VGND VPWR VPWR _17587_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13064__B1 _13040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14799_ _18089_/A _14798_/Y _25083_/Q _14798_/A VGND VGND VPWR VPWR _14799_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22323__B1 _20609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19326_ _19032_/A VGND VGND VPWR VPWR _19326_/X sky130_fd_sc_hd__buf_2
X_16538_ _16536_/Y _16533_/X _16537_/X _16533_/X VGND VGND VPWR VPWR _16538_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21080__A _15792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19257_ _18914_/A _13761_/X _13744_/X _13770_/X VGND VGND VPWR VPWR _19258_/A sky130_fd_sc_hd__or4_4
X_16469_ _16540_/A VGND VGND VPWR VPWR _16469_/X sky130_fd_sc_hd__buf_2
XANTENNA__17179__A2_N _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18208_ _18102_/A _18208_/B _18208_/C VGND VGND VPWR VPWR _18208_/X sky130_fd_sc_hd__and3_4
X_19188_ _23836_/Q VGND VGND VPWR VPWR _19188_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18139_ _18107_/A _18139_/B _18139_/C VGND VGND VPWR VPWR _18139_/X sky130_fd_sc_hd__and3_4
XFILLER_172_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21150_ _21031_/X _21149_/X VGND VGND VPWR VPWR _21150_/Y sky130_fd_sc_hd__nor2_4
XFILLER_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_90_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _24794_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12809__A1_N _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20101_ _20100_/Y VGND VGND VPWR VPWR _20101_/X sky130_fd_sc_hd__buf_2
X_21081_ _21081_/A VGND VGND VPWR VPWR _21082_/A sky130_fd_sc_hd__buf_2
XANTENNA__19255__B1 _19254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14422__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20032_ _20031_/Y _20029_/X _20010_/X _20029_/X VGND VGND VPWR VPWR _20032_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15816__B1 _24848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24840_ _24883_/CLK _24840_/D HRESETn VGND VGND VPWR VPWR _24840_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15831__A3 _16245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21983_ _21660_/X _21970_/X _21974_/Y _13793_/D _21982_/X VGND VGND VPWR VPWR _21983_/X
+ sky130_fd_sc_hd__a32o_4
X_24771_ _24777_/CLK _24771_/D HRESETn VGND VGND VPWR VPWR _22871_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24755__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16349__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20934_ _13659_/C _20929_/X _20933_/Y VGND VGND VPWR VPWR _20934_/Y sky130_fd_sc_hd__a21oi_4
X_23722_ _23716_/CLK _23722_/D VGND VGND VPWR VPWR _23722_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20865_/A _20865_/B VGND VGND VPWR VPWR _20865_/X sky130_fd_sc_hd__or2_4
X_23653_ _23642_/CLK _19716_/X VGND VGND VPWR VPWR _13458_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21117__A1 _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22314__B1 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _22754_/A _22601_/X _22604_/C VGND VGND VPWR VPWR _22625_/C sky130_fd_sc_hd__and3_4
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23565_/CLK _19915_/X VGND VGND VPWR VPWR _23584_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_169_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ _20788_/X _20795_/Y _15592_/A _20792_/X VGND VGND VPWR VPWR _24037_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_169_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22535_ _22535_/A _22535_/B VGND VGND VPWR VPWR _22535_/Y sky130_fd_sc_hd__nor2_4
X_25323_ _25181_/CLK _13501_/X HRESETn VGND VGND VPWR VPWR _25323_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20876__B1 _20863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22466_ _16259_/Y _22462_/X _15108_/Y _22459_/X VGND VGND VPWR VPWR _22467_/B sky130_fd_sc_hd__o22a_4
X_25254_ _25200_/CLK _13882_/X HRESETn VGND VGND VPWR VPWR _22129_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15898__A3 _16238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21140__D _13822_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22814__A _24601_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21417_ _21398_/X _20165_/Y VGND VGND VPWR VPWR _21417_/X sky130_fd_sc_hd__or2_4
X_24205_ _23654_/CLK _24205_/D HRESETn VGND VGND VPWR VPWR _18357_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18297__A1 _21834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25185_ _25177_/CLK _25185_/D HRESETn VGND VGND VPWR VPWR _14309_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22397_ _21785_/X _22396_/X _21277_/A VGND VGND VPWR VPWR _22397_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22533__B _21604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ _12150_/A VGND VGND VPWR VPWR _12150_/Y sky130_fd_sc_hd__inv_2
X_24136_ _24160_/CLK _18817_/X HRESETn VGND VGND VPWR VPWR _24136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18616__A1_N _16606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21348_ _21348_/A _21348_/B VGND VGND VPWR VPWR _21348_/X sky130_fd_sc_hd__or2_4
XFILLER_162_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11956__A _11934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_118_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24476_/CLK sky130_fd_sc_hd__clkbuf_1
X_12081_ _16193_/A _12081_/B _12109_/C _12080_/X VGND VGND VPWR VPWR _12081_/X sky130_fd_sc_hd__or4_4
X_24067_ _24500_/CLK _24067_/D HRESETn VGND VGND VPWR VPWR _24067_/Q sky130_fd_sc_hd__dfrtp_4
X_21279_ _21262_/X _21277_/X _21278_/X VGND VGND VPWR VPWR _21279_/X sky130_fd_sc_hd__a21o_4
XANTENNA__16956__A2_N _24293_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23018_ _24440_/Q _22947_/X _23015_/X _23017_/X VGND VGND VPWR VPWR _23018_/X sky130_fd_sc_hd__a211o_4
XFILLER_238_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15840_ _12333_/Y _15838_/X _15629_/X _15838_/X VGND VGND VPWR VPWR _24832_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15771_ _12523_/Y _15768_/X _15632_/X _15768_/X VGND VGND VPWR VPWR _24866_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12983_ _12796_/Y _12986_/B VGND VGND VPWR VPWR _12983_/Y sky130_fd_sc_hd__nand2_4
X_24969_ _24966_/CLK _24969_/D HRESETn VGND VGND VPWR VPWR _13915_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12787__A _25392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17510_ _25535_/Q _17585_/D _11768_/Y _24322_/Q VGND VGND VPWR VPWR _17510_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14722_ _14721_/X _13769_/X _14721_/X _13769_/X VGND VGND VPWR VPWR _14722_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11934_ _11933_/X VGND VGND VPWR VPWR _11934_/X sky130_fd_sc_hd__buf_2
X_18490_ _18490_/A _18490_/B VGND VGND VPWR VPWR _18492_/B sky130_fd_sc_hd__or2_4
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16232__B1 _15972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17441_ _17426_/A VGND VGND VPWR VPWR _17441_/X sky130_fd_sc_hd__buf_2
XANTENNA__23380__A _21023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14653_ _13617_/Y _14652_/Y _18016_/A _14652_/Y VGND VGND VPWR VPWR _14653_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11865_ HWDATA[2] VGND VGND VPWR VPWR _11865_/X sky130_fd_sc_hd__buf_2
XFILLER_72_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21108__B2 _21747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _19548_/A VGND VGND VPWR VPWR _19595_/A sky130_fd_sc_hd__buf_2
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17372_ _17364_/B _17364_/C _17298_/A _17369_/B VGND VGND VPWR VPWR _17372_/X sky130_fd_sc_hd__a211o_4
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ _25543_/Q VGND VGND VPWR VPWR _11796_/Y sky130_fd_sc_hd__inv_2
X_14584_ _14583_/X _14564_/X _13778_/A VGND VGND VPWR VPWR _14584_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19111_ _23863_/Q VGND VGND VPWR VPWR _21626_/B sky130_fd_sc_hd__inv_2
XPHY_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16323_ _16322_/Y _16320_/X _15965_/X _16320_/X VGND VGND VPWR VPWR _24637_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20867__B1 _20863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13535_ _14310_/A VGND VGND VPWR VPWR _13535_/Y sky130_fd_sc_hd__inv_2
X_19042_ _19041_/Y _19037_/X _18991_/X _19037_/X VGND VGND VPWR VPWR _23888_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12953__C _12855_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16254_ _22557_/A VGND VGND VPWR VPWR _16254_/Y sky130_fd_sc_hd__inv_2
X_13466_ _13217_/X _13464_/X _13465_/X VGND VGND VPWR VPWR _13466_/X sky130_fd_sc_hd__and3_4
XANTENNA__22724__A _22724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15205_ _14902_/A _15204_/Y VGND VGND VPWR VPWR _15205_/X sky130_fd_sc_hd__or2_4
XANTENNA__25284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ _12191_/Y _12414_/X VGND VGND VPWR VPWR _12417_/X sky130_fd_sc_hd__or2_4
XFILLER_127_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16185_ _16185_/A _16180_/X _16182_/X _16184_/X VGND VGND VPWR VPWR _16185_/X sky130_fd_sc_hd__or4_4
XFILLER_126_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17818__A _17762_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13397_ _13257_/X _13397_/B VGND VGND VPWR VPWR _13397_/X sky130_fd_sc_hd__or2_4
XANTENNA__16299__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_14_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__25213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _15311_/A _15134_/Y _24986_/Q _15135_/Y VGND VGND VPWR VPWR _15136_/X sky130_fd_sc_hd__a2bb2o_4
X_12348_ _12348_/A _12341_/X _12344_/X _12348_/D VGND VGND VPWR VPWR _12348_/X sky130_fd_sc_hd__or4_4
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_77_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23258__C _23253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11866__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _12278_/Y _22285_/A _12273_/X _21715_/A VGND VGND VPWR VPWR _12279_/X sky130_fd_sc_hd__a2bb2o_4
X_15067_ _15067_/A VGND VGND VPWR VPWR _15293_/A sky130_fd_sc_hd__buf_2
X_19944_ _19944_/A VGND VGND VPWR VPWR _22354_/B sky130_fd_sc_hd__inv_2
XANTENNA__14242__A _25202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12165__A1_N _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14018_ _14058_/C _14057_/A VGND VGND VPWR VPWR _14062_/C sky130_fd_sc_hd__or2_4
X_19875_ _19873_/Y _19874_/X _19807_/X _19874_/X VGND VGND VPWR VPWR _19875_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18826_ _18689_/C _18791_/B VGND VGND VPWR VPWR _18826_/Y sky130_fd_sc_hd__nand2_4
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16471__B1 _16385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18757_ _18776_/A _18757_/B _18756_/X VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__and3_4
XANTENNA__15813__A3 _15732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15969_ _12223_/Y _15962_/X _15967_/X _15968_/X VGND VGND VPWR VPWR _24772_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17708_ _17587_/Y _17610_/D _17611_/X _17705_/Y VGND VGND VPWR VPWR _17708_/X sky130_fd_sc_hd__a211o_4
XFILLER_36_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _24134_/Q VGND VGND VPWR VPWR _18689_/A sky130_fd_sc_hd__inv_2
XFILLER_224_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16223__B1 _15963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23290__A _23290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17639_ _17511_/A _17638_/Y VGND VGND VPWR VPWR _17639_/X sky130_fd_sc_hd__or2_4
XFILLER_210_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20650_ _20649_/X VGND VGND VPWR VPWR _20650_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15801__A _15826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19309_ _19301_/Y VGND VGND VPWR VPWR _19309_/X sky130_fd_sc_hd__buf_2
XFILLER_149_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20581_ _18883_/B _20579_/Y _20597_/C VGND VGND VPWR VPWR _20581_/X sky130_fd_sc_hd__and3_4
XFILLER_165_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22320_ _14441_/Y _22334_/B VGND VGND VPWR VPWR _22320_/Y sky130_fd_sc_hd__nor2_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22251_ _22266_/A _22246_/X _22250_/X VGND VGND VPWR VPWR _22251_/X sky130_fd_sc_hd__or3_4
XFILLER_191_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19476__B1 _19454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21202_ _21207_/A _19899_/Y VGND VGND VPWR VPWR _21204_/B sky130_fd_sc_hd__or2_4
X_22182_ _14487_/Y _14266_/A _25113_/Q _22190_/B VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11771__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21133_ _21119_/Y _21121_/X _21124_/X _21132_/X VGND VGND VPWR VPWR _21290_/A sky130_fd_sc_hd__a211o_4
XANTENNA__11776__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23024__A1 _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21064_ _21032_/X VGND VGND VPWR VPWR _21064_/X sky130_fd_sc_hd__buf_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20015_ _18290_/A _20015_/B _18283_/X _18294_/X VGND VGND VPWR VPWR _20016_/A sky130_fd_sc_hd__or4_4
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_28_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24823_ _24824_/CLK _24823_/D HRESETn VGND VGND VPWR VPWR _12613_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24754_ _24767_/CLK _15997_/X HRESETn VGND VGND VPWR VPWR _21451_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19400__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21966_ _22274_/A _21966_/B _21966_/C VGND VGND VPWR VPWR _21966_/X sky130_fd_sc_hd__or3_4
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _24206_/CLK _23705_/D VGND VGND VPWR VPWR _23705_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20900_/X _20916_/X _24502_/Q _20904_/X VGND VGND VPWR VPWR _20917_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _22228_/A _21894_/X _21896_/X VGND VGND VPWR VPWR _21897_/X sky130_fd_sc_hd__and3_4
X_24685_ _24684_/CLK _24685_/D HRESETn VGND VGND VPWR VPWR _13747_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15711__A _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _16720_/Y _20833_/X _20842_/X _20847_/X VGND VGND VPWR VPWR _20849_/A sky130_fd_sc_hd__o22a_4
X_23636_ _23916_/CLK _19767_/X VGND VGND VPWR VPWR _13179_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_230_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21432__B _21091_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20329__A _20323_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _13143_/C _13128_/X VGND VGND VPWR VPWR _20779_/X sky130_fd_sc_hd__or2_4
X_23567_ _24937_/CLK _23567_/D VGND VGND VPWR VPWR _19957_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13320_/A VGND VGND VPWR VPWR _13421_/A sky130_fd_sc_hd__buf_2
X_25306_ _25188_/CLK _25306_/D HRESETn VGND VGND VPWR VPWR _25306_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_155_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22518_ _16284_/X _22518_/B VGND VGND VPWR VPWR _22536_/A sky130_fd_sc_hd__nor2_4
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _23516_/CLK _20157_/X VGND VGND VPWR VPWR _20155_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22544__A _23148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13251_ _13468_/A _13251_/B VGND VGND VPWR VPWR _13251_/X sky130_fd_sc_hd__or2_4
X_22449_ _12778_/Y _22299_/B _22291_/B _12545_/Y _21431_/X VGND VGND VPWR VPWR _22449_/X
+ sky130_fd_sc_hd__o32a_4
X_25237_ _25246_/CLK _25237_/D HRESETn VGND VGND VPWR VPWR _14011_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__19467__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12202_ _22982_/A VGND VGND VPWR VPWR _12202_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13182_ _13182_/A VGND VGND VPWR VPWR _13416_/A sky130_fd_sc_hd__buf_2
X_25168_ _25168_/CLK _14359_/X HRESETn VGND VGND VPWR VPWR _14347_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12133_ _12132_/Y _12128_/X _11876_/X _12128_/X VGND VGND VPWR VPWR _25474_/D sky130_fd_sc_hd__a2bb2o_4
X_24119_ _24119_/CLK _20984_/X HRESETn VGND VGND VPWR VPWR _12160_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15158__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17990_ _17990_/A VGND VGND VPWR VPWR _18234_/A sky130_fd_sc_hd__buf_2
X_25099_ _25093_/CLK _14597_/X HRESETn VGND VGND VPWR VPWR _25099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12064_ _12108_/B VGND VGND VPWR VPWR _12081_/B sky130_fd_sc_hd__buf_2
X_16941_ _16941_/A _16941_/B _16939_/X _16940_/X VGND VGND VPWR VPWR _16941_/X sky130_fd_sc_hd__or4_4
XANTENNA__23375__A _23362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24677__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19660_ _19652_/Y VGND VGND VPWR VPWR _19660_/X sky130_fd_sc_hd__buf_2
X_16872_ _16866_/X VGND VGND VPWR VPWR _16872_/X sky130_fd_sc_hd__buf_2
XFILLER_237_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24606__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18611_ _16569_/Y _18737_/A _16569_/Y _18737_/A VGND VGND VPWR VPWR _18611_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16453__B1 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15823_ _12346_/Y _15821_/X _11797_/X _15821_/X VGND VGND VPWR VPWR _15823_/X sky130_fd_sc_hd__a2bb2o_4
X_19591_ _19591_/A VGND VGND VPWR VPWR _21194_/B sky130_fd_sc_hd__inv_2
X_18542_ _18471_/A _18540_/X _18541_/Y VGND VGND VPWR VPWR _24182_/D sky130_fd_sc_hd__o21a_4
XFILLER_218_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15754_ HWDATA[14] VGND VGND VPWR VPWR _15754_/X sky130_fd_sc_hd__buf_2
XFILLER_234_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12966_ _12777_/X _12952_/X _12891_/X _12962_/Y VGND VGND VPWR VPWR _12967_/A sky130_fd_sc_hd__a211o_4
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ _14728_/B VGND VGND VPWR VPWR _14707_/C sky130_fd_sc_hd__inv_2
X_11917_ _11890_/X _11887_/Y _11905_/X _17711_/B VGND VGND VPWR VPWR _11918_/A sky130_fd_sc_hd__a211o_4
X_18473_ _18534_/A _18531_/A _18472_/X VGND VGND VPWR VPWR _18473_/X sky130_fd_sc_hd__or3_4
XFILLER_206_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15685_ _15652_/Y _15678_/X _15656_/X _13680_/A _15684_/X VGND VGND VPWR VPWR _15685_/X
+ sky130_fd_sc_hd__a32o_4
X_12897_ _12780_/Y _12906_/B VGND VGND VPWR VPWR _12900_/B sky130_fd_sc_hd__or2_4
XFILLER_178_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17424_ _17424_/A VGND VGND VPWR VPWR _17424_/X sky130_fd_sc_hd__buf_2
XFILLER_233_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15621__A _15626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ _14635_/Y _13647_/X _25087_/Q _13645_/X VGND VGND VPWR VPWR _14637_/A sky130_fd_sc_hd__o22a_4
X_11848_ _11844_/Y _11845_/X _11847_/X _11845_/X VGND VGND VPWR VPWR _25531_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22157__C _22157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17252_/D _17355_/B VGND VGND VPWR VPWR _17391_/B sky130_fd_sc_hd__or2_4
X_14567_ _14567_/A VGND VGND VPWR VPWR _14593_/A sky130_fd_sc_hd__buf_2
X_11779_ _25548_/Q VGND VGND VPWR VPWR _11779_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16306_ HWDATA[26] VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__buf_2
X_13518_ _25315_/Q VGND VGND VPWR VPWR _13518_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17286_ _17203_/Y _17286_/B VGND VGND VPWR VPWR _17287_/C sky130_fd_sc_hd__or2_4
XFILLER_159_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14498_ _14496_/Y _14497_/X _14404_/X _14497_/X VGND VGND VPWR VPWR _14498_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19025_ _19024_/Y _19020_/X _18999_/X _19020_/A VGND VGND VPWR VPWR _19025_/X sky130_fd_sc_hd__a2bb2o_4
X_16237_ _22751_/A VGND VGND VPWR VPWR _16237_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13449_ _13417_/A _23933_/Q VGND VGND VPWR VPWR _13449_/X sky130_fd_sc_hd__or2_4
XFILLER_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20068__B2 _20065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16168_ _16166_/Y _16162_/X _15480_/X _16167_/X VGND VGND VPWR VPWR _16168_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11753__B1 _11752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15119_ _25010_/Q _24614_/Q _15318_/C _15118_/Y VGND VGND VPWR VPWR _15119_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15068__A _15293_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16099_ _16093_/Y _16098_/X _11752_/X _16098_/X VGND VGND VPWR VPWR _16099_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19927_ _19923_/Y _19926_/X _19790_/X _19926_/X VGND VGND VPWR VPWR _19927_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_101_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24824_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15218__D _15172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_164_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _24214_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17283__A _17243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19858_ _23604_/Q VGND VGND VPWR VPWR _19858_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16444__B1 _16073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18809_ _18809_/A _18809_/B VGND VGND VPWR VPWR _18810_/B sky130_fd_sc_hd__or2_4
XFILLER_84_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19789_ _19788_/Y VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__buf_2
XANTENNA__22517__B1 _15121_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21820_ _21493_/A _21818_/X _21820_/C VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__and3_4
XFILLER_237_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22629__A _22592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21751_ _16859_/Y _22146_/B _21591_/A _21750_/X VGND VGND VPWR VPWR _21751_/X sky130_fd_sc_hd__o22a_4
XFILLER_221_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20702_ _15645_/Y _20695_/X _20698_/X _20701_/Y VGND VGND VPWR VPWR _20702_/X sky130_fd_sc_hd__o22a_4
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21740__B2 _16731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21682_ _21682_/A _21682_/B VGND VGND VPWR VPWR _21682_/X sky130_fd_sc_hd__or2_4
X_24470_ _24430_/CLK _16763_/X HRESETn VGND VGND VPWR VPWR _24470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ _17399_/B _20632_/Y _20628_/X VGND VGND VPWR VPWR _20633_/X sky130_fd_sc_hd__and3_4
X_23421_ _24206_/CLK _20359_/X VGND VGND VPWR VPWR _23421_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19938__A _19925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23352_ _13811_/Y _14683_/A _13815_/Y _25062_/Q VGND VGND VPWR VPWR _23353_/A sky130_fd_sc_hd__o22a_4
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13981__A1 scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20564_ _14116_/A VGND VGND VPWR VPWR _20564_/X sky130_fd_sc_hd__buf_2
XFILLER_109_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22364__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22303_ _21314_/A VGND VGND VPWR VPWR _22303_/X sky130_fd_sc_hd__buf_2
XFILLER_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23283_ _21456_/X _23281_/X _22702_/X _23282_/X VGND VGND VPWR VPWR _23283_/X sky130_fd_sc_hd__o22a_4
XFILLER_153_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19449__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17458__A _24328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20495_ _20524_/A _23976_/D _20494_/Y VGND VGND VPWR VPWR _20520_/A sky130_fd_sc_hd__o21a_4
X_22234_ _14766_/X _20216_/Y VGND VGND VPWR VPWR _22234_/X sky130_fd_sc_hd__or2_4
X_25022_ _25018_/CLK _25022_/D HRESETn VGND VGND VPWR VPWR _15270_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_180_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22165_ _21116_/X _22158_/X _22161_/X _22164_/X VGND VGND VPWR VPWR _22165_/X sky130_fd_sc_hd__a211o_4
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_60_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21116_ _21872_/A VGND VGND VPWR VPWR _21116_/X sky130_fd_sc_hd__buf_2
XFILLER_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16683__B1 _16414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__A _21557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22096_ _21246_/A VGND VGND VPWR VPWR _22209_/A sky130_fd_sc_hd__buf_2
XANTENNA__24770__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22756__B1 _24875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21047_ _21046_/X VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__buf_2
XFILLER_59_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19621__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15789__A2 _15678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20782__A2 _20716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12820_ _12819_/Y _24807_/Q _12857_/A _12767_/Y VGND VGND VPWR VPWR _12824_/C sky130_fd_sc_hd__a2bb2o_4
X_24806_ _24794_/CLK _15897_/X HRESETn VGND VGND VPWR VPWR _24806_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13226__A _13423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22998_ _22732_/A VGND VGND VPWR VPWR _22998_/X sky130_fd_sc_hd__buf_2
XANTENNA__22539__A _23313_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12751_ _12955_/A VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__inv_2
X_24737_ _24738_/CLK _16045_/X HRESETn VGND VGND VPWR VPWR _16042_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21949_/A _21949_/B _21949_/C VGND VGND VPWR VPWR _21949_/X sky130_fd_sc_hd__and3_4
XFILLER_42_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16537__A _14427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11702_/A VGND VGND VPWR VPWR _13691_/A sky130_fd_sc_hd__inv_2
XFILLER_188_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _24963_/Q VGND VGND VPWR VPWR _15470_/Y sky130_fd_sc_hd__inv_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A VGND VGND VPWR VPWR _25426_/D sky130_fd_sc_hd__inv_2
X_24668_ _24666_/CLK _24668_/D HRESETn VGND VGND VPWR VPWR _24668_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14414_/Y _14418_/X _14420_/X _14418_/X VGND VGND VPWR VPWR _14421_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _23916_/CLK _23619_/D VGND VGND VPWR VPWR _19819_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_187_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24599_ _24601_/CLK _24599_/D HRESETn VGND VGND VPWR VPWR _16427_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _16969_/Y _17139_/X VGND VGND VPWR VPWR _17157_/A sky130_fd_sc_hd__or2_4
XFILLER_11_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14349_/C _14349_/D VGND VGND VPWR VPWR _14352_/X sky130_fd_sc_hd__or2_4
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22274__A _22274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13187_/X _13294_/X _13303_/C VGND VGND VPWR VPWR _13303_/X sky130_fd_sc_hd__and3_4
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ _16990_/A _17070_/Y VGND VGND VPWR VPWR _17073_/B sky130_fd_sc_hd__or2_4
X_14283_ _14282_/Y _14280_/X _14248_/X _14280_/X VGND VGND VPWR VPWR _25191_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16022_ _16021_/Y _16019_/X _11773_/X _16019_/X VGND VGND VPWR VPWR _24746_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13234_ _13228_/A VGND VGND VPWR VPWR _13356_/A sky130_fd_sc_hd__buf_2
XFILLER_108_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24858__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21798__B2 _22549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13165_ _13164_/Y VGND VGND VPWR VPWR _13451_/A sky130_fd_sc_hd__buf_2
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12305__A _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16674__B1 _16315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22721__B _22721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ _12123_/A VGND VGND VPWR VPWR _12116_/X sky130_fd_sc_hd__buf_2
X_13096_ _13002_/D _13102_/B VGND VGND VPWR VPWR _13096_/X sky130_fd_sc_hd__or2_4
X_17973_ _17973_/A VGND VGND VPWR VPWR _17973_/X sky130_fd_sc_hd__buf_2
X_12047_ _12047_/A VGND VGND VPWR VPWR _12047_/Y sky130_fd_sc_hd__inv_2
X_16924_ _22920_/A _24282_/Q _16127_/Y _16923_/Y VGND VGND VPWR VPWR _16924_/X sky130_fd_sc_hd__o22a_4
X_19712_ _19710_/Y _19711_/X _19566_/X _19711_/X VGND VGND VPWR VPWR _23655_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_237_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _23998_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16426__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20222__B2 _20219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16855_ _14954_/Y _16853_/X _16537_/X _16853_/X VGND VGND VPWR VPWR _16855_/X sky130_fd_sc_hd__a2bb2o_4
X_19643_ _19643_/A VGND VGND VPWR VPWR _19643_/X sky130_fd_sc_hd__buf_2
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15806_ _15826_/A VGND VGND VPWR VPWR _15806_/Y sky130_fd_sc_hd__inv_2
X_19574_ _19574_/A VGND VGND VPWR VPWR _19574_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14988__B1 _15258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16786_ _16785_/Y _16782_/X _16530_/X _16782_/X VGND VGND VPWR VPWR _16786_/X sky130_fd_sc_hd__a2bb2o_4
X_13998_ _25243_/Q VGND VGND VPWR VPWR _13998_/X sky130_fd_sc_hd__buf_2
XFILLER_93_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18525_ _18486_/D _18503_/X _18486_/B VGND VGND VPWR VPWR _18525_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21353__A _21353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15737_ _15758_/A VGND VGND VPWR VPWR _15737_/X sky130_fd_sc_hd__buf_2
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12949_ _12770_/Y _12609_/X VGND VGND VPWR VPWR _12988_/B sky130_fd_sc_hd__or2_4
XFILLER_34_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21722__B2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22168__B _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18456_ _18452_/X _18453_/X _18456_/C _18455_/X VGND VGND VPWR VPWR _18456_/X sky130_fd_sc_hd__or4_4
X_15668_ _15651_/X _15668_/B VGND VGND VPWR VPWR _15668_/X sky130_fd_sc_hd__or2_4
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17407_ _17407_/A _17407_/B VGND VGND VPWR VPWR _17408_/B sky130_fd_sc_hd__or2_4
X_14619_ _13561_/A _13593_/A VGND VGND VPWR VPWR _14619_/X sky130_fd_sc_hd__or2_4
X_18387_ _18386_/Y _18384_/X _24199_/Q _18384_/X VGND VGND VPWR VPWR _24200_/D sky130_fd_sc_hd__a2bb2o_4
X_15599_ _15599_/A VGND VGND VPWR VPWR _22934_/A sky130_fd_sc_hd__inv_2
X_17338_ _17338_/A _17317_/C VGND VGND VPWR VPWR _17341_/B sky130_fd_sc_hd__or2_4
XANTENNA__20289__B2 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21486__B1 _18306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17269_ _17345_/A _17277_/A VGND VGND VPWR VPWR _17283_/B sky130_fd_sc_hd__or2_4
X_19008_ _19148_/A VGND VGND VPWR VPWR _19008_/X sky130_fd_sc_hd__buf_2
X_20280_ _22385_/B _20279_/X _16866_/X _20279_/X VGND VGND VPWR VPWR _20280_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24599__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16910__A _16910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22631__B _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_47_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16665__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21528__A _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15526__A _15544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23970_ _23970_/CLK _23970_/D HRESETn VGND VGND VPWR VPWR _23970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22921_ _15800_/A _22920_/X _22503_/X _25544_/Q _22793_/X VGND VGND VPWR VPWR _22921_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22852_ _22941_/A VGND VGND VPWR VPWR _22852_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21803_ _21466_/X _21803_/B VGND VGND VPWR VPWR _21803_/X sky130_fd_sc_hd__or2_4
XANTENNA__21263__A _21263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22783_ _24806_/Q _22985_/B VGND VGND VPWR VPWR _22783_/X sky130_fd_sc_hd__or2_4
X_24522_ _24528_/CLK _24522_/D HRESETn VGND VGND VPWR VPWR _16627_/A sky130_fd_sc_hd__dfrtp_4
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21734_ _25252_/Q VGND VGND VPWR VPWR _21734_/Y sky130_fd_sc_hd__inv_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24453_ _24613_/CLK _16798_/X HRESETn VGND VGND VPWR VPWR _15019_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_169_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21665_ _21466_/X _21665_/B VGND VGND VPWR VPWR _21665_/X sky130_fd_sc_hd__or2_4
XANTENNA__12206__B2 _21091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23404_ _24217_/CLK _23404_/D VGND VGND VPWR VPWR _23404_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20616_ _20611_/X _20615_/X _20549_/B VGND VGND VPWR VPWR _20616_/X sky130_fd_sc_hd__o21a_4
X_21596_ _21596_/A _21596_/B VGND VGND VPWR VPWR _21610_/C sky130_fd_sc_hd__nor2_4
X_24384_ _24383_/CLK _24384_/D HRESETn VGND VGND VPWR VPWR _24384_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12109__B _12107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20547_ _14465_/A _23939_/Q VGND VGND VPWR VPWR _23935_/D sky130_fd_sc_hd__and2_4
X_23335_ _24515_/Q _16552_/A VGND VGND VPWR VPWR _23335_/Y sky130_fd_sc_hd__nor2_4
X_20478_ _20455_/C _20478_/B VGND VGND VPWR VPWR _20478_/X sky130_fd_sc_hd__or2_4
X_23266_ _16010_/A _21039_/X _21042_/X _23265_/X VGND VGND VPWR VPWR _23266_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16850__A1_N _14943_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25005_ _25002_/CLK _25005_/D HRESETn VGND VGND VPWR VPWR _25005_/Q sky130_fd_sc_hd__dfrtp_4
X_22217_ _21260_/A _22217_/B _22216_/X VGND VGND VPWR VPWR _22221_/B sky130_fd_sc_hd__and3_4
XFILLER_193_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23197_ _23113_/X _23196_/X _23159_/X _24852_/Q _23115_/X VGND VGND VPWR VPWR _23197_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22441__A2 _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16820__A _16810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16656__B1 _16294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22148_ _21607_/X _22146_/X _22148_/C VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__and3_4
XFILLER_160_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11964__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14970_ _14969_/Y VGND VGND VPWR VPWR _15243_/A sky130_fd_sc_hd__buf_2
X_22079_ _22380_/A _22077_/X _22078_/X VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__and3_4
XANTENNA__16865__A1_N _16864_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21157__B _21375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16408__B1 _16407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14682__A2 _13610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13921_ _13927_/A _13907_/Y _13917_/X _13927_/C _13920_/X VGND VGND VPWR VPWR _13921_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_48_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16640_ _16640_/A _16643_/A _16643_/B VGND VGND VPWR VPWR _16640_/X sky130_fd_sc_hd__or3_4
X_13852_ _13848_/A VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_67_0_HCLK clkbuf_8_66_0_HCLK/A VGND VGND VPWR VPWR _25443_/CLK sky130_fd_sc_hd__clkbuf_1
X_12803_ _12819_/A _12801_/Y _12952_/C _22139_/A VGND VGND VPWR VPWR _12803_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21173__A _15388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16571_ _16571_/A VGND VGND VPWR VPWR _16571_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13783_ _13607_/B VGND VGND VPWR VPWR _13828_/C sky130_fd_sc_hd__inv_2
XANTENNA__23091__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ _21675_/A _18310_/B VGND VGND VPWR VPWR _18310_/X sky130_fd_sc_hd__and2_4
X_15522_ _24943_/Q VGND VGND VPWR VPWR _15522_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _12713_/X _12734_/B _12741_/C VGND VGND VPWR VPWR _12734_/X sky130_fd_sc_hd__and3_4
X_19290_ _23800_/Q VGND VGND VPWR VPWR _21770_/B sky130_fd_sc_hd__inv_2
XFILLER_187_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18241_ _18248_/A VGND VGND VPWR VPWR _18241_/Y sky130_fd_sc_hd__inv_2
X_15453_ _15443_/A VGND VGND VPWR VPWR _15453_/X sky130_fd_sc_hd__buf_2
X_12665_ _12616_/B _12669_/B VGND VGND VPWR VPWR _12665_/Y sky130_fd_sc_hd__nand2_4
XFILLER_231_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _15486_/A VGND VGND VPWR VPWR _14404_/X sky130_fd_sc_hd__buf_2
XFILLER_230_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22716__B _22316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18172_ _15703_/X _18156_/X _18171_/X _24250_/Q _18029_/X VGND VGND VPWR VPWR _18172_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15384_/A _15384_/B _15384_/C VGND VGND VPWR VPWR _24996_/D sky130_fd_sc_hd__and3_4
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _25426_/Q VGND VGND VPWR VPWR _12596_/Y sky130_fd_sc_hd__inv_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ _24393_/Q _17122_/Y VGND VGND VPWR VPWR _17123_/X sky130_fd_sc_hd__or2_4
X_14335_ _25174_/Q _12172_/X _14334_/X VGND VGND VPWR VPWR _14335_/X sky130_fd_sc_hd__a21o_4
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23209__B2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17054_ _17047_/X _17054_/B _17054_/C VGND VGND VPWR VPWR _17055_/C sky130_fd_sc_hd__or3_4
XFILLER_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14266_ _14266_/A VGND VGND VPWR VPWR _21726_/B sky130_fd_sc_hd__buf_2
XANTENNA__24692__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16005_ _16004_/X VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__buf_2
X_13217_ _13164_/Y VGND VGND VPWR VPWR _13217_/X sky130_fd_sc_hd__buf_2
XANTENNA__24621__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14197_ _12061_/A _15558_/B VGND VGND VPWR VPWR _16378_/D sky130_fd_sc_hd__or2_4
XANTENNA__19833__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13148_ _20693_/B VGND VGND VPWR VPWR _20696_/B sky130_fd_sc_hd__inv_2
XANTENNA__21348__A _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11874__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13079_ _13051_/A VGND VGND VPWR VPWR _13104_/A sky130_fd_sc_hd__buf_2
X_17956_ _17944_/A _17956_/B VGND VGND VPWR VPWR _17956_/X sky130_fd_sc_hd__or2_4
XFILLER_239_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12133__B1 _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16907_ _17760_/C VGND VGND VPWR VPWR _17861_/C sky130_fd_sc_hd__buf_2
X_17887_ _16936_/X _17858_/B VGND VGND VPWR VPWR _17891_/B sky130_fd_sc_hd__or2_4
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19626_ _19626_/A VGND VGND VPWR VPWR _19626_/X sky130_fd_sc_hd__buf_2
XFILLER_238_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16838_ _24433_/Q VGND VGND VPWR VPWR _16838_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21083__A _21083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16769_ _15012_/Y _16768_/X _15748_/X _16768_/X VGND VGND VPWR VPWR _24467_/D sky130_fd_sc_hd__a2bb2o_4
X_19557_ _19565_/A VGND VGND VPWR VPWR _19557_/X sky130_fd_sc_hd__buf_2
XFILLER_207_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18508_ _18510_/B VGND VGND VPWR VPWR _18513_/B sky130_fd_sc_hd__inv_2
X_19488_ _19488_/A VGND VGND VPWR VPWR _22038_/B sky130_fd_sc_hd__inv_2
XFILLER_61_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21171__A2 _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18439_ _16244_/Y _18474_/A _16244_/Y _18474_/A VGND VGND VPWR VPWR _18443_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22626__B _22589_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21450_ _21311_/A VGND VGND VPWR VPWR _21450_/X sky130_fd_sc_hd__buf_2
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20401_ _21490_/B _20398_/X _19646_/A _20398_/X VGND VGND VPWR VPWR _20401_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21381_ _19617_/A _21971_/B _19568_/Y _21971_/B VGND VGND VPWR VPWR _21381_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24709__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14425__A _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20332_ _21953_/B _20329_/X _20000_/X _20329_/X VGND VGND VPWR VPWR _20332_/X sky130_fd_sc_hd__a2bb2o_4
X_23120_ _21436_/X VGND VGND VPWR VPWR _23120_/X sky130_fd_sc_hd__buf_2
XFILLER_190_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23051_ _23117_/A _23050_/X VGND VGND VPWR VPWR _23065_/B sky130_fd_sc_hd__and2_4
X_20263_ _20270_/A VGND VGND VPWR VPWR _20263_/X sky130_fd_sc_hd__buf_2
XFILLER_190_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22002_ _21853_/X _21880_/X _21893_/X _22002_/D VGND VGND VPWR VPWR HRDATA[4] sky130_fd_sc_hd__or4_4
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21631__B1 _14758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22974__A3 _22861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20194_ _20190_/Y _20193_/X _20102_/X _20193_/X VGND VGND VPWR VPWR _20194_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25172__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12124__B1 _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14664__A2 _14650_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23953_ _23954_/CLK _23953_/D HRESETn VGND VGND VPWR VPWR _20570_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_220_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _24613_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_244_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22904_ _16764_/A _22543_/A _22903_/X VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23884_ _23885_/CLK _23884_/D VGND VGND VPWR VPWR _23884_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22835_ _24738_/Q _21067_/X _21068_/X _22834_/X VGND VGND VPWR VPWR _22835_/X sky130_fd_sc_hd__a211o_4
XFILLER_213_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13504__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21698__B1 _21697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25554_ _25539_/CLK _25554_/D HRESETn VGND VGND VPWR VPWR _25554_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ _16691_/Y _22578_/B VGND VGND VPWR VPWR _22766_/X sky130_fd_sc_hd__and2_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21162__A2 _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24505_ _24503_/CLK _24505_/D HRESETn VGND VGND VPWR VPWR _16677_/A sky130_fd_sc_hd__dfrtp_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21717_ _21717_/A VGND VGND VPWR VPWR _21717_/Y sky130_fd_sc_hd__inv_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25485_ _24112_/CLK _12098_/X HRESETn VGND VGND VPWR VPWR _12097_/A sky130_fd_sc_hd__dfrtp_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22697_ _22535_/B _22697_/B VGND VGND VPWR VPWR _22697_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16815__A _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12222_/Y _12449_/X _12403_/X VGND VGND VPWR VPWR _12450_/Y sky130_fd_sc_hd__a21oi_4
X_24436_ _24437_/CLK _24436_/D HRESETn VGND VGND VPWR VPWR _14950_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18733__C _18733_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21648_ _21648_/A _20117_/Y VGND VGND VPWR VPWR _21649_/C sky130_fd_sc_hd__or2_4
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12381_ _25343_/Q VGND VGND VPWR VPWR _12381_/Y sky130_fd_sc_hd__inv_2
X_24367_ _24346_/CLK _24367_/D HRESETn VGND VGND VPWR VPWR _17186_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21579_ _12106_/A VGND VGND VPWR VPWR _21579_/X sky130_fd_sc_hd__buf_2
X_14120_ _14117_/X VGND VGND VPWR VPWR _14120_/X sky130_fd_sc_hd__buf_2
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23318_ _23299_/X _23302_/X _23306_/Y _23317_/X VGND VGND VPWR VPWR HRDATA[30] sky130_fd_sc_hd__a211o_4
XFILLER_153_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24298_ _25528_/CLK _17704_/X HRESETn VGND VGND VPWR VPWR _24298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22552__A _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17548__A1_N _11782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14051_ _25247_/Q _14015_/B _13999_/D _14014_/A VGND VGND VPWR VPWR _14052_/A sky130_fd_sc_hd__or4_4
X_23249_ _23249_/A _23248_/X VGND VGND VPWR VPWR _23258_/B sky130_fd_sc_hd__nor2_4
X_13002_ _12387_/X _12342_/Y _13002_/C _13002_/D VGND VGND VPWR VPWR _13002_/X sky130_fd_sc_hd__or4_4
XFILLER_180_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21168__A _18515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19291__B2 _19286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17810_ _17810_/A VGND VGND VPWR VPWR _17810_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18790_ _18687_/D _18733_/C VGND VGND VPWR VPWR _18791_/B sky130_fd_sc_hd__or2_4
X_17741_ _18290_/A _17733_/X _24224_/Q _17734_/Y VGND VGND VPWR VPWR _17741_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23383__A _21026_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14953_ _24420_/Q VGND VGND VPWR VPWR _14953_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13904_ _13936_/C VGND VGND VPWR VPWR _13923_/A sky130_fd_sc_hd__buf_2
XFILLER_247_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17381__A _24351_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17672_ _17701_/A _17529_/Y _17537_/Y _17671_/X VGND VGND VPWR VPWR _17672_/X sky130_fd_sc_hd__or4_4
X_14884_ _14883_/X VGND VGND VPWR VPWR _25048_/D sky130_fd_sc_hd__inv_2
X_16623_ _16623_/A VGND VGND VPWR VPWR _16623_/X sky130_fd_sc_hd__buf_2
X_19411_ _19409_/Y _19405_/X _19410_/X _19391_/X VGND VGND VPWR VPWR _23757_/D sky130_fd_sc_hd__a2bb2o_4
X_13835_ _13578_/Y _13831_/X _11818_/X _13834_/X VGND VGND VPWR VPWR _13835_/X sky130_fd_sc_hd__a2bb2o_4
X_16554_ _16554_/A VGND VGND VPWR VPWR _16554_/X sky130_fd_sc_hd__buf_2
X_19342_ _19340_/Y _19338_/X _19341_/X _19338_/X VGND VGND VPWR VPWR _19342_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ _13766_/A _25282_/Q VGND VGND VPWR VPWR _13767_/B sky130_fd_sc_hd__and2_4
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23301__A1_N _17270_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15505_ _16378_/A _15503_/X HADDR[21] _15503_/X VGND VGND VPWR VPWR _15505_/X sky130_fd_sc_hd__a2bb2o_4
X_12717_ _12621_/A _12723_/B VGND VGND VPWR VPWR _12718_/B sky130_fd_sc_hd__or2_4
X_19273_ _23806_/Q VGND VGND VPWR VPWR _21391_/B sky130_fd_sc_hd__inv_2
X_16485_ _24577_/Q VGND VGND VPWR VPWR _16485_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20361__B1 _15656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13697_ _13697_/A _13697_/B VGND VGND VPWR VPWR _13698_/B sky130_fd_sc_hd__or2_4
XFILLER_204_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16725__A _24485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18224_ _18060_/A _18224_/B VGND VGND VPWR VPWR _18226_/B sky130_fd_sc_hd__or2_4
X_15436_ _15436_/A VGND VGND VPWR VPWR _15436_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12648_ _12640_/B VGND VGND VPWR VPWR _12657_/A sky130_fd_sc_hd__buf_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24873__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18155_ _18059_/A _18151_/X _18154_/X VGND VGND VPWR VPWR _18155_/X sky130_fd_sc_hd__or3_4
XFILLER_178_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11869__A _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15367_ _15362_/A _15361_/X _15324_/X _15363_/Y VGND VGND VPWR VPWR _15367_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24802__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12579_ _25419_/Q VGND VGND VPWR VPWR _12579_/Y sky130_fd_sc_hd__inv_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18940__A _18952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17106_ _17106_/A _17104_/X _17106_/C VGND VGND VPWR VPWR _24399_/D sky130_fd_sc_hd__and3_4
X_14318_ _14315_/X _14317_/Y _25329_/Q _14315_/X VGND VGND VPWR VPWR _25183_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18086_ _18191_/A _18083_/X _18086_/C VGND VGND VPWR VPWR _18087_/C sky130_fd_sc_hd__and3_4
X_15298_ _15387_/A VGND VGND VPWR VPWR _15355_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_112_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17037_ _24403_/Q VGND VGND VPWR VPWR _17037_/Y sky130_fd_sc_hd__inv_2
X_14249_ _14247_/Y _14245_/X _14248_/X _14245_/X VGND VGND VPWR VPWR _14249_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23277__B _23274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18988_ _23905_/Q VGND VGND VPWR VPWR _18988_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21806__A _21668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17939_ _18023_/A _23892_/Q VGND VGND VPWR VPWR _17939_/X sky130_fd_sc_hd__or2_4
XFILLER_239_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13854__B1 _13812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17291__A _17345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15804__A _15796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20950_ _20947_/Y _20948_/Y _20949_/X VGND VGND VPWR VPWR _20950_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19609_ _21971_/A _19606_/X _19560_/X _19606_/X VGND VGND VPWR VPWR _19609_/X sky130_fd_sc_hd__a2bb2o_4
X_20881_ _20881_/A VGND VGND VPWR VPWR _20904_/A sky130_fd_sc_hd__inv_2
XFILLER_242_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_50_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _24233_/CLK sky130_fd_sc_hd__clkbuf_1
X_22620_ _22620_/A VGND VGND VPWR VPWR _22620_/Y sky130_fd_sc_hd__inv_2
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21541__A _15792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22551_ _21288_/X _22549_/X _21968_/X _22550_/X VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__o22a_4
XFILLER_195_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21502_ _21497_/A _21502_/B VGND VGND VPWR VPWR _21502_/X sky130_fd_sc_hd__or2_4
XANTENNA__19011__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25270_ _25281_/CLK _25270_/D HRESETn VGND VGND VPWR VPWR _25270_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22482_ _21090_/A VGND VGND VPWR VPWR _23322_/B sky130_fd_sc_hd__buf_2
XFILLER_194_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24221_ _24295_/CLK _18296_/X HRESETn VGND VGND VPWR VPWR _24221_/Q sky130_fd_sc_hd__dfrtp_4
X_21433_ _22202_/C VGND VGND VPWR VPWR _22986_/A sky130_fd_sc_hd__buf_2
XANTENNA__21447__A3 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21364_ _18393_/Y _21580_/A _12175_/A _12106_/A VGND VGND VPWR VPWR _21364_/X sky130_fd_sc_hd__o22a_4
X_24152_ _24966_/CLK _18757_/X HRESETn VGND VGND VPWR VPWR _24152_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21852__B1 _21565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20315_ _20302_/Y VGND VGND VPWR VPWR _20315_/X sky130_fd_sc_hd__buf_2
X_23103_ _21879_/A _23100_/X _23102_/X VGND VGND VPWR VPWR _23103_/X sky130_fd_sc_hd__and3_4
XFILLER_174_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15531__B1 HADDR[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21295_ _21295_/A VGND VGND VPWR VPWR _21322_/A sky130_fd_sc_hd__inv_2
X_24083_ _25543_/CLK _20479_/X HRESETn VGND VGND VPWR VPWR _13782_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16370__A _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20246_ _20245_/Y _20240_/X _19753_/X _20240_/X VGND VGND VPWR VPWR _23464_/D sky130_fd_sc_hd__a2bb2o_4
X_23034_ _21427_/A _23032_/Y _22844_/X _23033_/X VGND VGND VPWR VPWR _23035_/A sky130_fd_sc_hd__o22a_4
XFILLER_162_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _20172_/A VGND VGND VPWR VPWR _20177_/X sky130_fd_sc_hd__buf_2
XFILLER_131_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15834__A1 _15833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15834__B2 _15802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19025__B2 _19020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24985_ _24975_/CLK _15422_/Y HRESETn VGND VGND VPWR VPWR _15153_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13845__B1 _13844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15714__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ _20003_/A VGND VGND VPWR VPWR _19639_/A sky130_fd_sc_hd__buf_2
X_23936_ _24012_/CLK _23936_/D HRESETn VGND VGND VPWR VPWR _22115_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15598__B1 _11790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _11880_/Y VGND VGND VPWR VPWR _11881_/X sky130_fd_sc_hd__buf_2
X_23867_ _23628_/CLK _23867_/D VGND VGND VPWR VPWR _19102_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_189_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13620_ _18098_/A VGND VGND VPWR VPWR _18023_/A sky130_fd_sc_hd__buf_2
XFILLER_244_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13234__A _13228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22818_ _24435_/Q _21085_/A _22815_/X _22817_/X VGND VGND VPWR VPWR _22818_/X sky130_fd_sc_hd__a211o_4
X_23798_ _23926_/CLK _23798_/D VGND VGND VPWR VPWR _23798_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_198_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13551_ _24258_/Q _13550_/X VGND VGND VPWR VPWR _13551_/X sky130_fd_sc_hd__and2_4
X_25537_ _24386_/CLK _25537_/D HRESETn VGND VGND VPWR VPWR _11820_/A sky130_fd_sc_hd__dfrtp_4
X_22749_ _22527_/X _22746_/X _22431_/X _22748_/X VGND VGND VPWR VPWR _22750_/A sky130_fd_sc_hd__o22a_4
XFILLER_186_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12502_ _12502_/A VGND VGND VPWR VPWR _12503_/B sky130_fd_sc_hd__inv_2
X_16270_ _16268_/Y _16264_/X _15480_/X _16269_/X VGND VGND VPWR VPWR _24656_/D sky130_fd_sc_hd__a2bb2o_4
X_13482_ _13474_/Y _13480_/Y _13481_/X _13480_/Y VGND VGND VPWR VPWR _25330_/D sky130_fd_sc_hd__a2bb2o_4
X_25468_ _25456_/CLK _12405_/Y HRESETn VGND VGND VPWR VPWR _25468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15221_ _15075_/D _15220_/X VGND VGND VPWR VPWR _15221_/X sky130_fd_sc_hd__or2_4
X_12433_ _25461_/Q _12432_/Y VGND VGND VPWR VPWR _12433_/X sky130_fd_sc_hd__or2_4
X_24419_ _24613_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _24419_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15770__B1 _15629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25399_ _25402_/CLK _25399_/D HRESETn VGND VGND VPWR VPWR _25399_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15152_ _15345_/C _15158_/A _24991_/Q _15095_/Y VGND VGND VPWR VPWR _15152_/X sky130_fd_sc_hd__a2bb2o_4
X_12364_ _13038_/A _24848_/Q _13038_/A _24848_/Q VGND VGND VPWR VPWR _12369_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23378__A _23378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22282__A _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14103_ _14103_/A VGND VGND VPWR VPWR _14116_/A sky130_fd_sc_hd__inv_2
XFILLER_154_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22713__C _21752_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15083_ _15082_/Y _16434_/A _15082_/Y _16434_/A VGND VGND VPWR VPWR _15091_/A sky130_fd_sc_hd__a2bb2o_4
X_19960_ _19960_/A VGND VGND VPWR VPWR _19960_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _12208_/Y _12255_/Y _12222_/Y _12197_/A VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__or4_4
XFILLER_153_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14034_ _14062_/A _14031_/Y _14054_/C _14034_/D VGND VGND VPWR VPWR _14034_/X sky130_fd_sc_hd__or4_4
X_18911_ _18910_/Y _18907_/X _17452_/X _18907_/X VGND VGND VPWR VPWR _23933_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19891_ _21937_/B _19888_/X _19636_/X _19888_/X VGND VGND VPWR VPWR _23593_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12823__A2_N _22755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18842_ _16474_/A _24160_/Q _16474_/Y _18720_/A VGND VGND VPWR VPWR _18842_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15985_ _12230_/Y _15983_/X _15765_/X _15983_/X VGND VGND VPWR VPWR _24762_/D sky130_fd_sc_hd__a2bb2o_4
X_18773_ _18773_/A VGND VGND VPWR VPWR _18773_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13836__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14936_ _14936_/A VGND VGND VPWR VPWR _14936_/Y sky130_fd_sc_hd__inv_2
X_17724_ _24217_/Q VGND VGND VPWR VPWR _21210_/A sky130_fd_sc_hd__buf_2
XFILLER_36_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12838__A2_N _21712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18000__A _18008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ _14823_/A _14823_/B _14823_/A _14823_/B VGND VGND VPWR VPWR _14868_/A sky130_fd_sc_hd__a2bb2o_4
X_17655_ _17646_/C _17646_/D VGND VGND VPWR VPWR _17656_/C sky130_fd_sc_hd__nand2_4
XFILLER_208_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_37_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_74_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13818_ _13818_/A VGND VGND VPWR VPWR _16729_/A sky130_fd_sc_hd__buf_2
X_16606_ _16606_/A VGND VGND VPWR VPWR _16606_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17586_ _24300_/Q VGND VGND VPWR VPWR _17588_/B sky130_fd_sc_hd__inv_2
X_14798_ _14798_/A VGND VGND VPWR VPWR _14798_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22457__A _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16537_ _14427_/A VGND VGND VPWR VPWR _16537_/X sky130_fd_sc_hd__buf_2
X_19325_ _19324_/Y VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__buf_2
X_13749_ _13749_/A VGND VGND VPWR VPWR _13749_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22176__B _22176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16468_ _16468_/A _16468_/B VGND VGND VPWR VPWR _16540_/A sky130_fd_sc_hd__nor2_4
X_19256_ _23812_/Q VGND VGND VPWR VPWR _22372_/B sky130_fd_sc_hd__inv_2
XFILLER_188_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15419_ _24986_/Q _15419_/B VGND VGND VPWR VPWR _15420_/B sky130_fd_sc_hd__or2_4
X_18207_ _18013_/A _18207_/B VGND VGND VPWR VPWR _18208_/C sky130_fd_sc_hd__or2_4
XFILLER_148_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19187_ _19186_/Y _19181_/X _19139_/X _19181_/A VGND VGND VPWR VPWR _23837_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19766__A _19765_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16399_ _16397_/Y _16398_/X _16306_/X _16398_/X VGND VGND VPWR VPWR _24611_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18138_ _18138_/A _18138_/B _18137_/X VGND VGND VPWR VPWR _18139_/C sky130_fd_sc_hd__or3_4
XFILLER_145_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18069_ _18069_/A _18069_/B _18068_/X VGND VGND VPWR VPWR _18069_/X sky130_fd_sc_hd__and3_4
X_20100_ _13764_/X VGND VGND VPWR VPWR _20100_/Y sky130_fd_sc_hd__inv_2
X_21080_ _15792_/X VGND VGND VPWR VPWR _21081_/A sky130_fd_sc_hd__inv_2
XFILLER_171_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20031_ _20031_/A VGND VGND VPWR VPWR _20031_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13319__A _13356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12223__A _22910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24770_ _24777_/CLK _15973_/X HRESETn VGND VGND VPWR VPWR _24770_/Q sky130_fd_sc_hd__dfrtp_4
X_21982_ _21978_/Y _21979_/X _21980_/X _21981_/X VGND VGND VPWR VPWR _21982_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23173__D _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _23716_/CLK _23721_/D VGND VGND VPWR VPWR _23721_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ _20907_/B _20933_/B VGND VGND VPWR VPWR _20933_/Y sky130_fd_sc_hd__nor2_4
XFILLER_215_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23916_/CLK _23652_/D VGND VGND VPWR VPWR _13173_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _20865_/A VGND VGND VPWR VPWR _20864_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24795__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21117__A2 _21113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18518__B1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22314__A1 _16615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22603_ _16603_/A _23303_/B _21755_/A _22602_/X VGND VGND VPWR VPWR _22604_/C sky130_fd_sc_hd__a211o_4
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _23582_/CLK _23583_/D VGND VGND VPWR VPWR _23583_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_223_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22865__A2 _22531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24724__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20795_ _13129_/C _20790_/X _20794_/Y VGND VGND VPWR VPWR _20795_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16365__A _16290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25322_ _25177_/CLK _13503_/X HRESETn VGND VGND VPWR VPWR _13502_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_168_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22534_ _22534_/A VGND VGND VPWR VPWR _22535_/B sky130_fd_sc_hd__buf_2
XFILLER_179_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25253_ _25253_/CLK _13884_/X HRESETn VGND VGND VPWR VPWR _21847_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19676__A _19675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22465_ _21596_/A _22464_/X VGND VGND VPWR VPWR _22465_/Y sky130_fd_sc_hd__nor2_4
XFILLER_148_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24204_ _23654_/CLK _18375_/X HRESETn VGND VGND VPWR VPWR _18372_/A sky130_fd_sc_hd__dfrtp_4
X_21416_ _21412_/A _21414_/X _21415_/X VGND VGND VPWR VPWR _21416_/X sky130_fd_sc_hd__and3_4
X_25184_ _25177_/CLK _14313_/Y HRESETn VGND VGND VPWR VPWR _25184_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22396_ _22373_/A _22392_/X _22393_/X _22394_/X _22395_/X VGND VGND VPWR VPWR _22396_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20189__A2_N _20184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24135_ _24160_/CLK _18819_/Y HRESETn VGND VGND VPWR VPWR _24135_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15504__B1 HADDR[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21347_ _16460_/A _21340_/X _21347_/C VGND VGND VPWR VPWR _21425_/B sky130_fd_sc_hd__and3_4
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12080_ _12080_/A VGND VGND VPWR VPWR _12080_/X sky130_fd_sc_hd__buf_2
X_24066_ _24500_/CLK _24066_/D HRESETn VGND VGND VPWR VPWR _13658_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21278_ _17455_/X VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__buf_2
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22830__A _24569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23017_ _24472_/Q _23016_/X _22903_/X VGND VGND VPWR VPWR _23017_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20229_ _21394_/B _20226_/X _19810_/A _20226_/X VGND VGND VPWR VPWR _23470_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15770_ _12551_/Y _15768_/X _15629_/X _15768_/X VGND VGND VPWR VPWR _24867_/D sky130_fd_sc_hd__a2bb2o_4
X_12982_ _12837_/Y _12984_/B _12981_/Y VGND VGND VPWR VPWR _12982_/X sky130_fd_sc_hd__o21a_4
X_24968_ _24975_/CLK _24968_/D HRESETn VGND VGND VPWR VPWR _13955_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14491__B1 _14427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14721_ _22214_/A VGND VGND VPWR VPWR _14721_/X sky130_fd_sc_hd__buf_2
XFILLER_218_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22553__B2 _21322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11933_ _11933_/A _11908_/Y VGND VGND VPWR VPWR _11933_/X sky130_fd_sc_hd__and2_4
X_23919_ _23918_/CLK _18953_/X VGND VGND VPWR VPWR _23919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24899_ _24015_/CLK _24899_/D HRESETn VGND VGND VPWR VPWR _15645_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_217_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ _17440_/A VGND VGND VPWR VPWR _21567_/A sky130_fd_sc_hd__inv_2
XFILLER_217_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14652_ _14650_/C VGND VGND VPWR VPWR _14652_/Y sky130_fd_sc_hd__inv_2
X_11864_ _25527_/Q VGND VGND VPWR VPWR _11864_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14243__B1 _13809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13603_/A _13603_/B VGND VGND VPWR VPWR _19548_/A sky130_fd_sc_hd__or2_4
X_17371_ _17363_/A _17371_/B _17370_/X VGND VGND VPWR VPWR _17371_/X sky130_fd_sc_hd__and3_4
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _14593_/A _14582_/Y _14586_/C _25102_/Q VGND VGND VPWR VPWR _14583_/X sky130_fd_sc_hd__and4_4
XFILLER_186_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ _11792_/Y _11786_/X _11793_/X _11794_/X VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15991__B1 _15636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19182__B1 _19091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ _16322_/A VGND VGND VPWR VPWR _16322_/Y sky130_fd_sc_hd__inv_2
X_19110_ _21771_/B _19105_/X _16890_/X _19105_/X VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ _25311_/Q _20972_/B _13533_/X VGND VGND VPWR VPWR _25311_/D sky130_fd_sc_hd__a21o_4
XFILLER_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19041_ _18125_/B VGND VGND VPWR VPWR _19041_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16253_ _16250_/Y _16251_/X _16252_/X _16251_/X VGND VGND VPWR VPWR _24663_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13465_ _13245_/X _13465_/B VGND VGND VPWR VPWR _13465_/X sky130_fd_sc_hd__or2_4
XANTENNA__15743__B1 _11790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15204_ _15203_/X VGND VGND VPWR VPWR _15204_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22724__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12416_ _12191_/A _12415_/Y VGND VGND VPWR VPWR _12418_/B sky130_fd_sc_hd__or2_4
XANTENNA__21816__B1 _18306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16184_ _13599_/B _16184_/B VGND VGND VPWR VPWR _16184_/X sky130_fd_sc_hd__and2_4
X_13396_ _13249_/A _13396_/B VGND VGND VPWR VPWR _13398_/B sky130_fd_sc_hd__or2_4
XFILLER_127_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15135_ _15135_/A VGND VGND VPWR VPWR _15135_/Y sky130_fd_sc_hd__inv_2
X_12347_ _25358_/Q _24843_/Q _13068_/A _12346_/Y VGND VGND VPWR VPWR _12348_/D sky130_fd_sc_hd__o22a_4
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15066_ _15065_/X VGND VGND VPWR VPWR _25045_/D sky130_fd_sc_hd__inv_2
X_19943_ _19942_/Y _19938_/X _19856_/X _19925_/Y VGND VGND VPWR VPWR _23573_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12278_ _25444_/Q VGND VGND VPWR VPWR _12278_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22740__A _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ _14021_/B _13998_/X _14000_/C _14022_/A VGND VGND VPWR VPWR _14057_/A sky130_fd_sc_hd__or4_4
XFILLER_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22241__B1 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _19861_/Y VGND VGND VPWR VPWR _19874_/X sky130_fd_sc_hd__buf_2
XFILLER_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18825_ _18806_/A _18825_/B _18824_/Y VGND VGND VPWR VPWR _24133_/D sky130_fd_sc_hd__and3_4
XFILLER_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21356__A _14229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _18756_/A _18756_/B VGND VGND VPWR VPWR _18756_/X sky130_fd_sc_hd__or2_4
X_15968_ _15947_/A VGND VGND VPWR VPWR _15968_/X sky130_fd_sc_hd__buf_2
X_17707_ _17703_/B _17706_/X _17702_/C VGND VGND VPWR VPWR _17707_/X sky130_fd_sc_hd__and3_4
X_14919_ _14919_/A _14911_/X _14915_/X _14918_/X VGND VGND VPWR VPWR _14919_/X sky130_fd_sc_hd__or4_4
X_15899_ _15894_/X _15895_/X _16241_/A _22726_/A _15896_/X VGND VGND VPWR VPWR _15899_/X
+ sky130_fd_sc_hd__a32o_4
X_18687_ _18797_/A _18648_/A _18685_/Y _18687_/D VGND VGND VPWR VPWR _18687_/X sky130_fd_sc_hd__or4_4
X_17638_ _17637_/X VGND VGND VPWR VPWR _17638_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14234__B1 _13844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21091__A _21091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17569_ _17569_/A _17569_/B VGND VGND VPWR VPWR _17569_/X sky130_fd_sc_hd__or2_4
XFILLER_210_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19308_ _19151_/A VGND VGND VPWR VPWR _19308_/X sky130_fd_sc_hd__buf_2
XFILLER_177_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20580_ _18891_/X VGND VGND VPWR VPWR _20597_/C sky130_fd_sc_hd__buf_2
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_124_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _24473_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_220_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_187_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _24121_/CLK sky130_fd_sc_hd__clkbuf_1
X_19239_ _19238_/Y _19236_/X _19148_/X _19236_/X VGND VGND VPWR VPWR _23819_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20820__A1_N _20698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12218__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22250_ _22265_/A _22247_/X _22250_/C VGND VGND VPWR VPWR _22250_/X sky130_fd_sc_hd__and3_4
XFILLER_191_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21201_ _17714_/A _21199_/X _21200_/X VGND VGND VPWR VPWR _21201_/X sky130_fd_sc_hd__and3_4
X_22181_ _22181_/A VGND VGND VPWR VPWR _22181_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21132_ _21605_/A _21126_/X _21132_/C VGND VGND VPWR VPWR _21132_/X sky130_fd_sc_hd__and3_4
XFILLER_132_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23024__A2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21063_ _21063_/A VGND VGND VPWR VPWR _21079_/A sky130_fd_sc_hd__buf_2
XFILLER_235_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13049__A _13049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20014_ _23548_/Q VGND VGND VPWR VPWR _22351_/B sky130_fd_sc_hd__inv_2
XFILLER_113_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18987__B1 _17433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12888__A _12888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11792__A _25544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24822_ _24824_/CLK _15857_/X HRESETn VGND VGND VPWR VPWR _12989_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_228_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14473__B1 _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24753_ _24757_/CLK _24753_/D HRESETn VGND VGND VPWR VPWR _21091_/A sky130_fd_sc_hd__dfrtp_4
X_21965_ _21961_/X _21964_/X _18306_/A VGND VGND VPWR VPWR _21966_/C sky130_fd_sc_hd__o21a_4
XANTENNA__24905__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23704_ _23703_/CLK _23704_/D VGND VGND VPWR VPWR _23704_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20914_/Y _20911_/X _20915_/X VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__o21a_4
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24684_ _24684_/CLK _16188_/X HRESETn VGND VGND VPWR VPWR _14769_/A sky130_fd_sc_hd__dfrtp_4
X_21896_ _21895_/X _21896_/B VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__or2_4
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16511__A1_N _16510_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_20_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23644_/CLK _19770_/X VGND VGND VPWR VPWR _13260_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20846_/Y _13662_/X _13664_/X VGND VGND VPWR VPWR _20847_/X sky130_fd_sc_hd__o21a_4
XFILLER_199_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15973__B1 _15972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19164__B1 _19139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_83_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23566_ _24937_/CLK _19961_/X VGND VGND VPWR VPWR _19960_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_195_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20778_ _20761_/X _20777_/X _15601_/A _20765_/X VGND VGND VPWR VPWR _20778_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18911__B1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25305_ _23615_/CLK _13656_/X HRESETn VGND VGND VPWR VPWR _25305_/Q sky130_fd_sc_hd__dfrtp_4
X_22517_ _16256_/Y _22462_/A _15121_/Y _22459_/A VGND VGND VPWR VPWR _22518_/B sky130_fd_sc_hd__o22a_4
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23513_/CLK _23497_/D VGND VGND VPWR VPWR _23497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16526__A1_N _16524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23983__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ _13443_/A VGND VGND VPWR VPWR _13468_/A sky130_fd_sc_hd__buf_2
X_25236_ _25105_/CLK _25236_/D HRESETn VGND VGND VPWR VPWR _14011_/A sky130_fd_sc_hd__dfrtp_4
X_22448_ _12213_/Y _22425_/B _22284_/X _12327_/Y _21547_/X VGND VGND VPWR VPWR _22448_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_183_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12201_ _25448_/Q _12199_/Y _12299_/A _24779_/Q VGND VGND VPWR VPWR _12207_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13181_ _13200_/A _13179_/X _13181_/C VGND VGND VPWR VPWR _13181_/X sky130_fd_sc_hd__and3_4
X_25167_ _24121_/CLK _14362_/Y HRESETn VGND VGND VPWR VPWR _25167_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22471__B1 _13822_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22379_ _22095_/A _22379_/B VGND VGND VPWR VPWR _22379_/X sky130_fd_sc_hd__or2_4
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _12132_/A VGND VGND VPWR VPWR _12132_/Y sky130_fd_sc_hd__inv_2
X_24118_ _24119_/CLK _20983_/X HRESETn VGND VGND VPWR VPWR _24118_/Q sky130_fd_sc_hd__dfrtp_4
X_25098_ _25093_/CLK _14600_/X HRESETn VGND VGND VPWR VPWR _25098_/Q sky130_fd_sc_hd__dfrtp_4
X_12063_ _21583_/B VGND VGND VPWR VPWR _12108_/B sky130_fd_sc_hd__buf_2
X_16940_ _16140_/Y _24277_/Q _16140_/Y _24277_/Q VGND VGND VPWR VPWR _16940_/X sky130_fd_sc_hd__a2bb2o_4
X_24049_ _24488_/CLK _20845_/Y HRESETn VGND VGND VPWR VPWR _13660_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18978__B1 _18908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16871_ _16870_/X VGND VGND VPWR VPWR _16871_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18610_ _18681_/A VGND VGND VPWR VPWR _18737_/A sky130_fd_sc_hd__buf_2
XFILLER_219_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15822_ _12324_/Y _15818_/X _11793_/X _15821_/X VGND VGND VPWR VPWR _15822_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16453__B2 _16384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19590_ _21505_/B _19587_/X _11964_/X _19587_/X VGND VGND VPWR VPWR _19590_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14464__B1 _14420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15753_ _15737_/X _15751_/X _15752_/X _24875_/Q _15749_/X VGND VGND VPWR VPWR _15753_/X
+ sky130_fd_sc_hd__a32o_4
X_18541_ _18471_/A _18540_/X _18494_/X VGND VGND VPWR VPWR _18541_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21904__A _22093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12965_ _12984_/A _12963_/X _12964_/X VGND VGND VPWR VPWR _12965_/X sky130_fd_sc_hd__and3_4
XANTENNA__24646__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11916_ _11881_/X _11914_/X _11905_/X _11913_/Y VGND VGND VPWR VPWR _25520_/D sky130_fd_sc_hd__a2bb2o_4
X_14704_ _21630_/A _14703_/X _21630_/A _14703_/X VGND VGND VPWR VPWR _14728_/B sky130_fd_sc_hd__a2bb2o_4
X_15684_ _15651_/X _15683_/X VGND VGND VPWR VPWR _15684_/X sky130_fd_sc_hd__or2_4
X_18472_ _18540_/A _18540_/B _18472_/C VGND VGND VPWR VPWR _18472_/X sky130_fd_sc_hd__or3_4
XFILLER_73_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12896_ _12817_/Y _12895_/X VGND VGND VPWR VPWR _12906_/B sky130_fd_sc_hd__or2_4
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14635_ _25087_/Q VGND VGND VPWR VPWR _14635_/Y sky130_fd_sc_hd__inv_2
X_17423_ _21373_/A VGND VGND VPWR VPWR _17424_/A sky130_fd_sc_hd__buf_2
X_11847_ _11847_/A VGND VGND VPWR VPWR _11847_/X sky130_fd_sc_hd__buf_2
XANTENNA__15964__B1 _15963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25149__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14595_/A VGND VGND VPWR VPWR _14566_/X sky130_fd_sc_hd__buf_2
X_17354_ _17193_/Y VGND VGND VPWR VPWR _17364_/B sky130_fd_sc_hd__buf_2
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11775_/Y _11769_/X _11776_/X _11777_/X VGND VGND VPWR VPWR _25549_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13517_ _12009_/Y _13516_/X _11856_/X _13516_/X VGND VGND VPWR VPWR _25316_/D sky130_fd_sc_hd__a2bb2o_4
X_16305_ _16325_/A VGND VGND VPWR VPWR _16305_/X sky130_fd_sc_hd__buf_2
X_17285_ _24375_/Q _17284_/Y VGND VGND VPWR VPWR _17285_/X sky130_fd_sc_hd__or2_4
X_14497_ _14485_/A VGND VGND VPWR VPWR _14497_/X sky130_fd_sc_hd__buf_2
XANTENNA__16733__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16236_ _16233_/Y _16235_/X _11805_/X _16235_/X VGND VGND VPWR VPWR _24668_/D sky130_fd_sc_hd__a2bb2o_4
X_19024_ _19024_/A VGND VGND VPWR VPWR _19024_/Y sky130_fd_sc_hd__inv_2
X_13448_ _13416_/A _13448_/B _13447_/X VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__or3_4
XFILLER_174_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16167_ _16096_/X VGND VGND VPWR VPWR _16167_/X sky130_fd_sc_hd__buf_2
XANTENNA__25434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ _13411_/A _23855_/Q VGND VGND VPWR VPWR _13379_/X sky130_fd_sc_hd__or2_4
XFILLER_126_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15118_ _24614_/Q VGND VGND VPWR VPWR _15118_/Y sky130_fd_sc_hd__inv_2
X_16098_ _16097_/X VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__buf_2
XANTENNA__21017__A1 _23980_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15049_ _15043_/X _15044_/X _15049_/C _15049_/D VGND VGND VPWR VPWR _15064_/B sky130_fd_sc_hd__or4_4
X_19926_ _19925_/Y VGND VGND VPWR VPWR _19926_/X sky130_fd_sc_hd__buf_2
XFILLER_123_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21086__A _21172_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19857_ _21241_/B _19851_/X _19856_/X _19838_/Y VGND VGND VPWR VPWR _23605_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18808_ _18808_/A VGND VGND VPWR VPWR _24139_/D sky130_fd_sc_hd__inv_2
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19788_ _19788_/A VGND VGND VPWR VPWR _19788_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21814__A _21676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18739_ _18739_/A _18739_/B _18739_/C VGND VGND VPWR VPWR _24156_/D sky130_fd_sc_hd__and3_4
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12858__D _12834_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21750_ _16794_/Y _21589_/B VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__and2_4
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20701_ _13131_/A _13131_/B _13132_/B VGND VGND VPWR VPWR _20701_/Y sky130_fd_sc_hd__a21oi_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21681_ _21936_/A VGND VGND VPWR VPWR _21682_/A sky130_fd_sc_hd__buf_2
XFILLER_224_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15955__B1 _24779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14428__A _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12769__B1 _12888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13570__A1_N _25265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23420_ _24206_/CLK _23420_/D VGND VGND VPWR VPWR _20360_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_211_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13332__A _13423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20632_ _17398_/A _17398_/B VGND VGND VPWR VPWR _20632_/Y sky130_fd_sc_hd__nand2_4
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23351_ _14561_/X _23351_/B VGND VGND VPWR VPWR _24079_/D sky130_fd_sc_hd__or2_4
XFILLER_220_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20563_ _20563_/A VGND VGND VPWR VPWR _23951_/D sky130_fd_sc_hd__inv_2
XFILLER_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22302_ _22302_/A _21091_/B VGND VGND VPWR VPWR _22302_/X sky130_fd_sc_hd__or2_4
X_23282_ _16102_/Y _22569_/X _22861_/X _11757_/Y _22864_/X VGND VGND VPWR VPWR _23282_/X
+ sky130_fd_sc_hd__o32a_4
X_20494_ _24010_/Q VGND VGND VPWR VPWR _20494_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25021_ _25018_/CLK _15274_/Y HRESETn VGND VGND VPWR VPWR _14924_/A sky130_fd_sc_hd__dfrtp_4
X_22233_ _22226_/A _22233_/B VGND VGND VPWR VPWR _22235_/B sky130_fd_sc_hd__or2_4
XANTENNA__11787__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22164_ _21063_/A _22163_/X VGND VGND VPWR VPWR _22164_/X sky130_fd_sc_hd__and2_4
XFILLER_105_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21115_ _21321_/A VGND VGND VPWR VPWR _21872_/A sky130_fd_sc_hd__inv_2
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22095_ _22095_/A _20197_/Y VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__or2_4
XFILLER_114_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21708__B _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22756__A1 _21058_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22756__B2 _22565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21046_ _21046_/A VGND VGND VPWR VPWR _21046_/X sky130_fd_sc_hd__buf_2
XFILLER_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15789__A3 _15782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22508__B2 _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24805_ _24794_/CLK _24805_/D HRESETn VGND VGND VPWR VPWR _22755_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_234_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21724__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22997_ _23208_/A _22984_/X _22997_/C _22996_/X VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__or4_4
XFILLER_243_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15534__A2_N _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12750_ _21023_/A _12403_/X _12749_/Y VGND VGND VPWR VPWR _12750_/X sky130_fd_sc_hd__o21a_4
X_24736_ _24738_/CLK _16047_/X HRESETn VGND VGND VPWR VPWR _24736_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15722__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21948_ _21948_/A _19953_/Y VGND VGND VPWR VPWR _21949_/C sky130_fd_sc_hd__or2_4
XANTENNA__24057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _13698_/A _22525_/A _13698_/A _22525_/A VGND VGND VPWR VPWR _11708_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12596_/Y _12676_/B _12657_/A _12678_/B VGND VGND VPWR VPWR _12682_/A sky130_fd_sc_hd__a211o_4
X_24667_ _24666_/CLK _24667_/D HRESETn VGND VGND VPWR VPWR _22751_/A sky130_fd_sc_hd__dfrtp_4
X_21879_ _21879_/A _21879_/B _21878_/X VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__and3_4
XFILLER_70_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14338__A _14338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19137__B1 _19048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A VGND VGND VPWR VPWR _14420_/X sky130_fd_sc_hd__buf_2
XANTENNA__13242__A _13153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _25507_/CLK _23618_/D VGND VGND VPWR VPWR _19821_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12224__A2 _22910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24598_ _24601_/CLK _16431_/X HRESETn VGND VGND VPWR VPWR _16430_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22287__A3 _21308_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _12169_/D _14350_/Y _14359_/A VGND VGND VPWR VPWR _25170_/D sky130_fd_sc_hd__o21a_4
XFILLER_156_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23549_ _24217_/CLK _23549_/D VGND VGND VPWR VPWR _20012_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22692__B1 _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13171_/X _13298_/X _13301_/X VGND VGND VPWR VPWR _13303_/C sky130_fd_sc_hd__or3_4
X_17070_ _17072_/B VGND VGND VPWR VPWR _17070_/Y sky130_fd_sc_hd__inv_2
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _25191_/Q VGND VGND VPWR VPWR _14282_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_170_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24100_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16371__B1 _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16021_ _16021_/A VGND VGND VPWR VPWR _16021_/Y sky130_fd_sc_hd__inv_2
X_13233_ _13153_/X VGND VGND VPWR VPWR _13322_/A sky130_fd_sc_hd__buf_2
X_25219_ _23395_/CLK _25219_/D HRESETn VGND VGND VPWR VPWR _25219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_27_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _25528_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12179__A1_N _12168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ _13211_/A VGND VGND VPWR VPWR _13164_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22290__A _21719_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12115_ _25481_/Q VGND VGND VPWR VPWR _12140_/A sky130_fd_sc_hd__inv_2
XANTENNA__22721__C _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ _12339_/Y _13104_/B VGND VGND VPWR VPWR _13102_/B sky130_fd_sc_hd__or2_4
X_17972_ _17954_/X _17969_/X _18031_/A _24254_/Q _17973_/A VGND VGND VPWR VPWR _17972_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24898__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19711_ _19698_/Y VGND VGND VPWR VPWR _19711_/X sky130_fd_sc_hd__buf_2
XFILLER_111_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22747__B2 _21322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12046_ _12045_/Y _12043_/X _12047_/A _12043_/X VGND VGND VPWR VPWR _12046_/X sky130_fd_sc_hd__a2bb2o_4
X_16923_ _24282_/Q VGND VGND VPWR VPWR _16923_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24827__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19642_ _19624_/Y VGND VGND VPWR VPWR _19642_/X sky130_fd_sc_hd__buf_2
XFILLER_93_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16854_ _14899_/Y _16853_/X _16534_/X _16853_/X VGND VGND VPWR VPWR _16854_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15805_ _15790_/X _15804_/X _15723_/X _24855_/Q _15802_/X VGND VGND VPWR VPWR _24855_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21634__A _22388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19573_ _18282_/X _19480_/X _19505_/X VGND VGND VPWR VPWR _19574_/A sky130_fd_sc_hd__or3_4
XANTENNA__24480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ _14012_/A VGND VGND VPWR VPWR _14032_/A sky130_fd_sc_hd__buf_2
X_16785_ _24458_/Q VGND VGND VPWR VPWR _16785_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14988__B2 _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18524_ _18492_/A _18517_/B _18524_/C VGND VGND VPWR VPWR _18524_/X sky130_fd_sc_hd__and3_4
XANTENNA__15632__A _14423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12948_ _12988_/A VGND VGND VPWR VPWR _12984_/A sky130_fd_sc_hd__buf_2
X_15736_ _12548_/Y _15730_/X _11776_/X _15730_/X VGND VGND VPWR VPWR _15736_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18455_ _16263_/Y _24169_/Q _16271_/Y _24166_/Q VGND VGND VPWR VPWR _18455_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12879_ _12878_/X VGND VGND VPWR VPWR _12880_/B sky130_fd_sc_hd__inv_2
X_15667_ _15667_/A VGND VGND VPWR VPWR _15668_/B sky130_fd_sc_hd__buf_2
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14248__A _14248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _20668_/A _17406_/B VGND VGND VPWR VPWR _17407_/B sky130_fd_sc_hd__or2_4
X_14618_ _14571_/B _14617_/Y _14566_/X _14611_/X _13575_/A VGND VGND VPWR VPWR _25090_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_178_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15598_ _15596_/Y _15597_/X _11790_/X _15597_/X VGND VGND VPWR VPWR _24918_/D sky130_fd_sc_hd__a2bb2o_4
X_18386_ _18386_/A VGND VGND VPWR VPWR _18386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15070__C _15258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22465__A _21596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14549_ scl_oen_o_S4 _14543_/X _14544_/Y _14548_/Y VGND VGND VPWR VPWR _14550_/B
+ sky130_fd_sc_hd__o22a_4
X_17337_ _17336_/X VGND VGND VPWR VPWR _24362_/D sky130_fd_sc_hd__inv_2
XANTENNA__22683__B1 _21591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17268_ _17294_/A _17267_/X VGND VGND VPWR VPWR _17277_/A sky130_fd_sc_hd__or2_4
XANTENNA__16362__B1 _16073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17278__B _17243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19007_ HWDATA[6] VGND VGND VPWR VPWR _19148_/A sky130_fd_sc_hd__buf_2
X_16219_ _16219_/A VGND VGND VPWR VPWR _16219_/Y sky130_fd_sc_hd__inv_2
X_17199_ _24624_/Q _24353_/Q _16356_/Y _17198_/X VGND VGND VPWR VPWR _17200_/D sky130_fd_sc_hd__o22a_4
XFILLER_162_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16114__B1 _11773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17294__A _17294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21528__B _21425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19909_ _19909_/A VGND VGND VPWR VPWR _19909_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24568__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22920_ _22920_/A _22882_/X VGND VGND VPWR VPWR _22920_/X sky130_fd_sc_hd__or2_4
XFILLER_229_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21544__A _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22851_ _11747_/A VGND VGND VPWR VPWR _22851_/X sky130_fd_sc_hd__buf_2
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21802_ _21795_/Y _21801_/Y _13804_/C VGND VGND VPWR VPWR _21841_/C sky130_fd_sc_hd__o21a_4
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22782_ _22306_/A VGND VGND VPWR VPWR _23056_/A sky130_fd_sc_hd__buf_2
XANTENNA__21174__B1 _21332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21713__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24521_ _24556_/CLK _16630_/X HRESETn VGND VGND VPWR VPWR _24521_/Q sky130_fd_sc_hd__dfrtp_4
X_21733_ _21733_/A _21733_/B VGND VGND VPWR VPWR _21733_/Y sky130_fd_sc_hd__nor2_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20921__B1 _20863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24452_ _24613_/CLK _16800_/X HRESETn VGND VGND VPWR VPWR _24452_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21664_ _21652_/Y _21663_/Y _13804_/C VGND VGND VPWR VPWR _21708_/C sky130_fd_sc_hd__o21a_4
X_23403_ _23400_/CLK _23403_/D VGND VGND VPWR VPWR _22408_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_138_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20615_ _20609_/A _20612_/Y _20613_/Y _14504_/X _20614_/X VGND VGND VPWR VPWR _20615_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24383_ _24383_/CLK _24383_/D HRESETn VGND VGND VPWR VPWR _17159_/A sky130_fd_sc_hd__dfrtp_4
X_21595_ _22459_/A _21590_/X _22462_/A _21594_/X VGND VGND VPWR VPWR _21596_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23334_ _12188_/A _21082_/X _23332_/X _23333_/X _22510_/C VGND VGND VPWR VPWR _23334_/X
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__11965__B2 _11934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20546_ _24095_/Q _20451_/X _20515_/X VGND VGND VPWR VPWR _20546_/X sky130_fd_sc_hd__a21o_4
XFILLER_193_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16353__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_243_0_HCLK clkbuf_8_242_0_HCLK/A VGND VGND VPWR VPWR _23976_/CLK sky130_fd_sc_hd__clkbuf_1
X_23265_ _16296_/A _22954_/B _22830_/C VGND VGND VPWR VPWR _23265_/X sky130_fd_sc_hd__and3_4
X_20477_ _20477_/A _20461_/C _20477_/C VGND VGND VPWR VPWR _20478_/B sky130_fd_sc_hd__and3_4
XFILLER_192_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25004_ _25002_/CLK _25004_/D HRESETn VGND VGND VPWR VPWR _15354_/A sky130_fd_sc_hd__dfrtp_4
X_22216_ _21259_/A _19928_/Y VGND VGND VPWR VPWR _22216_/X sky130_fd_sc_hd__or2_4
XANTENNA__12531__A2_N _24876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16105__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21719__A _24620_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23196_ _23196_/A _22669_/B VGND VGND VPWR VPWR _23196_/X sky130_fd_sc_hd__or2_4
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22441__A3 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22147_ _22986_/A VGND VGND VPWR VPWR _22148_/C sky130_fd_sc_hd__buf_2
XANTENNA__15717__A _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22078_ _22095_/A _22078_/B VGND VGND VPWR VPWR _22078_/X sky130_fd_sc_hd__or2_4
XANTENNA__24920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13237__A _13282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13920_ _13923_/A _13927_/B _13927_/A _13907_/Y VGND VGND VPWR VPWR _13920_/X sky130_fd_sc_hd__o22a_4
X_21029_ _21029_/A VGND VGND VPWR VPWR _22306_/A sky130_fd_sc_hd__buf_2
XFILLER_247_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13851_ _13558_/Y _13848_/X _13806_/X _13848_/X VGND VGND VPWR VPWR _25264_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19358__B1 _19246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _25378_/Q VGND VGND VPWR VPWR _12952_/C sky130_fd_sc_hd__inv_2
X_13782_ _13782_/A VGND VGND VPWR VPWR _16464_/B sky130_fd_sc_hd__buf_2
X_16570_ _16569_/Y _16567_/X _16309_/X _16567_/X VGND VGND VPWR VPWR _24545_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21173__B _21173_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ _25411_/Q _12733_/B VGND VGND VPWR VPWR _12734_/B sky130_fd_sc_hd__or2_4
X_15521_ _15519_/Y _15520_/X HADDR[14] _15520_/X VGND VGND VPWR VPWR _15521_/X sky130_fd_sc_hd__a2bb2o_4
X_24719_ _24787_/CLK _24719_/D HRESETn VGND VGND VPWR VPWR _24719_/Q sky130_fd_sc_hd__dfrtp_4
X_15452_ _13951_/A _15446_/X _15441_/X _13934_/X _15447_/X VGND VGND VPWR VPWR _15452_/X
+ sky130_fd_sc_hd__a32o_4
X_18240_ _21974_/A _20405_/A VGND VGND VPWR VPWR _18248_/A sky130_fd_sc_hd__or2_4
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12664_ _12616_/A _12666_/B _12663_/Y VGND VGND VPWR VPWR _25431_/D sky130_fd_sc_hd__o21a_4
XFILLER_203_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14103_/A _14390_/B VGND VGND VPWR VPWR _14403_/X sky130_fd_sc_hd__or2_4
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_53_0_HCLK clkbuf_5_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _15383_/A _15383_/B VGND VGND VPWR VPWR _15384_/C sky130_fd_sc_hd__or2_4
X_18171_ _18107_/A _18163_/X _18171_/C VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__and3_4
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12595_/A VGND VGND VPWR VPWR _12595_/Y sky130_fd_sc_hd__inv_2
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _14334_/A VGND VGND VPWR VPWR _14334_/X sky130_fd_sc_hd__buf_2
X_17122_ _17110_/B VGND VGND VPWR VPWR _17122_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16344__B1 _16248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17053_ _17139_/A _17051_/Y _17053_/C _17052_/Y VGND VGND VPWR VPWR _17054_/C sky130_fd_sc_hd__or4_4
XFILLER_156_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14265_ _21375_/A VGND VGND VPWR VPWR _14266_/A sky130_fd_sc_hd__buf_2
XFILLER_171_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22417__B1 _22415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16004_ _16003_/X VGND VGND VPWR VPWR _16004_/X sky130_fd_sc_hd__buf_2
X_13216_ _13454_/A _13213_/X _13216_/C VGND VGND VPWR VPWR _13225_/B sky130_fd_sc_hd__and3_4
XFILLER_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14196_ _12061_/B VGND VGND VPWR VPWR _15558_/B sky130_fd_sc_hd__inv_2
XFILLER_152_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13147_ _13147_/A _13147_/B VGND VGND VPWR VPWR _20693_/B sky130_fd_sc_hd__or2_4
XANTENNA__21348__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18003__A _18234_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13078_ _13077_/X VGND VGND VPWR VPWR _13078_/Y sky130_fd_sc_hd__inv_2
X_17955_ _18023_/A _17955_/B VGND VGND VPWR VPWR _17955_/X sky130_fd_sc_hd__or2_4
XANTENNA__24661__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12029_ _12029_/A VGND VGND VPWR VPWR _12029_/Y sky130_fd_sc_hd__inv_2
X_16906_ _24273_/Q VGND VGND VPWR VPWR _17760_/C sky130_fd_sc_hd__inv_2
X_17886_ _17886_/A VGND VGND VPWR VPWR _24267_/D sky130_fd_sc_hd__inv_2
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19625_ _19624_/Y VGND VGND VPWR VPWR _19625_/X sky130_fd_sc_hd__buf_2
X_16837_ _16836_/Y _16834_/X _15752_/X _16834_/X VGND VGND VPWR VPWR _24434_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16458__A _16192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15083__B1 _15082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19349__B1 _19326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19556_ _23706_/Q VGND VGND VPWR VPWR _19556_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21083__B _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16768_ _16782_/A VGND VGND VPWR VPWR _16768_/X sky130_fd_sc_hd__buf_2
XFILLER_207_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18507_ _18507_/A VGND VGND VPWR VPWR _18507_/Y sky130_fd_sc_hd__inv_2
X_15719_ _15725_/A VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__buf_2
XFILLER_206_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19769__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19487_ _22244_/B _19484_/X _11943_/X _19484_/X VGND VGND VPWR VPWR _19487_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16699_ _16699_/A VGND VGND VPWR VPWR _16699_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18438_ _18432_/X _18435_/X _18436_/X _18438_/D VGND VGND VPWR VPWR _18438_/X sky130_fd_sc_hd__or4_4
XFILLER_22_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21459__A1 _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18369_ _18365_/Y _18368_/Y _18364_/X _18368_/A VGND VGND VPWR VPWR _24207_/D sky130_fd_sc_hd__o22a_4
XANTENNA__25205__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16193__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20400_ _20400_/A VGND VGND VPWR VPWR _21490_/B sky130_fd_sc_hd__inv_2
XFILLER_175_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21380_ _21380_/A VGND VGND VPWR VPWR _21971_/B sky130_fd_sc_hd__buf_2
XANTENNA__16335__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15138__B2 _16432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20331_ _20331_/A VGND VGND VPWR VPWR _21953_/B sky130_fd_sc_hd__inv_2
XFILLER_134_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16886__B2 _16877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23050_ _22777_/X _23049_/X _22872_/X _24848_/Q _22779_/X VGND VGND VPWR VPWR _23050_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_10_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23529_/CLK sky130_fd_sc_hd__clkbuf_1
X_20262_ _13275_/B VGND VGND VPWR VPWR _20262_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23081__B1 _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24749__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22001_ _22000_/X VGND VGND VPWR VPWR _22002_/D sky130_fd_sc_hd__inv_2
Xclkbuf_8_73_0_HCLK clkbuf_8_73_0_HCLK/A VGND VGND VPWR VPWR _24765_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15537__A _21135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20193_ _20193_/A VGND VGND VPWR VPWR _20193_/X sky130_fd_sc_hd__buf_2
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15256__B _15172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17752__A _17752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23952_ _23960_/CLK _23952_/D HRESETn VGND VGND VPWR VPWR _20566_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_243_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22903_ _21335_/X VGND VGND VPWR VPWR _22903_/X sky130_fd_sc_hd__buf_2
XFILLER_244_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18260__B1 _17433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23883_ _23880_/CLK _23883_/D VGND VGND VPWR VPWR _23883_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16368__A _14412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22834_ _24634_/Q _23027_/B _22513_/B VGND VGND VPWR VPWR _22834_/X sky130_fd_sc_hd__and3_4
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25553_ _24697_/CLK _11764_/X HRESETn VGND VGND VPWR VPWR _25553_/Q sky130_fd_sc_hd__dfrtp_4
X_22765_ _15608_/Y _22577_/B VGND VGND VPWR VPWR _22765_/X sky130_fd_sc_hd__and2_4
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24504_ _24500_/CLK _24504_/D HRESETn VGND VGND VPWR VPWR _24504_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21716_ _15565_/X _21715_/X _21445_/X _24828_/Q _21341_/X VGND VGND VPWR VPWR _21717_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25484_ _24112_/CLK _12100_/X HRESETn VGND VGND VPWR VPWR _12099_/A sky130_fd_sc_hd__dfrtp_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22696_ _21124_/X _22694_/X _21229_/X _22695_/X VGND VGND VPWR VPWR _22697_/B sky130_fd_sc_hd__o22a_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ _24431_/CLK _24435_/D HRESETn VGND VGND VPWR VPWR _24435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21647_ _21625_/A _21647_/B VGND VGND VPWR VPWR _21647_/X sky130_fd_sc_hd__or2_4
XFILLER_184_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12380_ _12380_/A _12374_/X _12380_/C _12380_/D VGND VGND VPWR VPWR _12380_/X sky130_fd_sc_hd__or4_4
X_24366_ _24346_/CLK _24366_/D HRESETn VGND VGND VPWR VPWR _17229_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16326__B1 _15967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21578_ _21577_/X VGND VGND VPWR VPWR _21578_/X sky130_fd_sc_hd__buf_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22833__A _17212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23317_ _23156_/A _23317_/B _23317_/C _23317_/D VGND VGND VPWR VPWR _23317_/X sky130_fd_sc_hd__or4_4
XFILLER_193_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20529_ _20473_/B _20528_/X _20513_/X VGND VGND VPWR VPWR _20529_/X sky130_fd_sc_hd__o21a_4
X_24297_ _24937_/CLK _17707_/X HRESETn VGND VGND VPWR VPWR _24297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14050_ _14050_/A VGND VGND VPWR VPWR _14554_/A sky130_fd_sc_hd__inv_2
X_23248_ _20818_/A _23006_/X _20956_/Y _22808_/X VGND VGND VPWR VPWR _23248_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17646__B _17578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13001_ _25350_/Q VGND VGND VPWR VPWR _13002_/D sky130_fd_sc_hd__inv_2
XFILLER_140_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23179_ _23137_/X _23177_/X _23139_/X _23178_/X VGND VGND VPWR VPWR _23180_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21168__B _21173_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19083__A2_N _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17740_ _17740_/A VGND VGND VPWR VPWR _18290_/A sky130_fd_sc_hd__buf_2
XANTENNA__17662__A _17691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14952_ _25030_/Q _14950_/Y _15275_/A _14954_/A VGND VGND VPWR VPWR _14960_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13903_ _13902_/X VGND VGND VPWR VPWR _13903_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17671_ _17567_/Y _17587_/Y VGND VGND VPWR VPWR _17671_/X sky130_fd_sc_hd__or2_4
XANTENNA__24001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14883_ _14877_/Y _14819_/X _14820_/X _14882_/X VGND VGND VPWR VPWR _14883_/X sky130_fd_sc_hd__o22a_4
X_19410_ _19139_/A VGND VGND VPWR VPWR _19410_/X sky130_fd_sc_hd__buf_2
X_16622_ _16622_/A VGND VGND VPWR VPWR _16622_/Y sky130_fd_sc_hd__inv_2
X_13834_ _13838_/A VGND VGND VPWR VPWR _13834_/X sky130_fd_sc_hd__buf_2
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19341_ _19048_/A VGND VGND VPWR VPWR _19341_/X sky130_fd_sc_hd__buf_2
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13765_ _19837_/A _13757_/X _13764_/X VGND VGND VPWR VPWR _13765_/Y sky130_fd_sc_hd__o21ai_4
X_16553_ _16623_/A VGND VGND VPWR VPWR _16554_/A sky130_fd_sc_hd__buf_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19751__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ _15558_/B _15500_/X HADDR[22] _15503_/X VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12716_ _12725_/A _12715_/X VGND VGND VPWR VPWR _12723_/B sky130_fd_sc_hd__or2_4
X_19272_ _19270_/Y _19271_/X _16894_/X _19271_/X VGND VGND VPWR VPWR _23807_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13696_ _11676_/Y _13695_/X VGND VGND VPWR VPWR _13697_/B sky130_fd_sc_hd__or2_4
X_16484_ _16482_/Y _16483_/X _16306_/X _16483_/X VGND VGND VPWR VPWR _16484_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16565__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18223_ _18191_/A _18223_/B _18222_/X VGND VGND VPWR VPWR _18227_/B sky130_fd_sc_hd__and3_4
XFILLER_176_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12647_ _12630_/A _12630_/B _12642_/B _12647_/D VGND VGND VPWR VPWR _12647_/X sky130_fd_sc_hd__or4_4
X_15435_ _13944_/A _15435_/B _13948_/C VGND VGND VPWR VPWR _15436_/A sky130_fd_sc_hd__or3_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15366_ _15384_/A _15364_/X _15366_/C VGND VGND VPWR VPWR _25002_/D sky130_fd_sc_hd__and3_4
X_18154_ _17975_/X _18152_/X _18154_/C VGND VGND VPWR VPWR _18154_/X sky130_fd_sc_hd__and3_4
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12578_ _12570_/X _12578_/B _12578_/C _12577_/X VGND VGND VPWR VPWR _12608_/A sky130_fd_sc_hd__or4_4
XFILLER_8_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22743__A _22592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20113__B2 _20109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _17105_/A _17102_/X VGND VGND VPWR VPWR _17106_/C sky130_fd_sc_hd__or2_4
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14317_ MSO_S2 _14316_/X _25182_/Q _14311_/X VGND VGND VPWR VPWR _14317_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15297_ _15293_/A _15256_/X _15297_/C VGND VGND VPWR VPWR _15297_/X sky130_fd_sc_hd__and3_4
X_18085_ _18084_/X _23905_/Q VGND VGND VPWR VPWR _18086_/C sky130_fd_sc_hd__or2_4
XFILLER_144_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14248_ _14248_/A VGND VGND VPWR VPWR _14248_/X sky130_fd_sc_hd__buf_2
X_17036_ _24401_/Q VGND VGND VPWR VPWR _17057_/A sky130_fd_sc_hd__inv_2
XANTENNA__24842__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _14174_/A VGND VGND VPWR VPWR _14179_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18987_ _18985_/Y _18986_/X _17433_/X _18986_/X VGND VGND VPWR VPWR _23906_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22169__A2 _21312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17938_ _13639_/X VGND VGND VPWR VPWR _17954_/A sky130_fd_sc_hd__buf_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17869_ _17861_/B _17861_/D VGND VGND VPWR VPWR _17872_/B sky130_fd_sc_hd__or2_4
XFILLER_238_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19608_ _19608_/A VGND VGND VPWR VPWR _21971_/A sky130_fd_sc_hd__inv_2
XFILLER_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20880_ _24057_/Q _13668_/X _20879_/Y VGND VGND VPWR VPWR _20880_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_199_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14803__B1 _25062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19539_ _21826_/B _19534_/X _11957_/X _19534_/X VGND VGND VPWR VPWR _19539_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22637__B _22589_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22550_ _22550_/A _22595_/B VGND VGND VPWR VPWR _22550_/X sky130_fd_sc_hd__and2_4
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21501_ _21466_/X _21501_/B VGND VGND VPWR VPWR _21501_/X sky130_fd_sc_hd__or2_4
X_22481_ _22452_/X _22458_/X _22465_/Y _22480_/X VGND VGND VPWR VPWR HRDATA[8] sky130_fd_sc_hd__a211o_4
XFILLER_195_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24220_ _23565_/CLK _24220_/D HRESETn VGND VGND VPWR VPWR _18319_/A sky130_fd_sc_hd__dfrtp_4
X_21432_ _21432_/A _21091_/B VGND VGND VPWR VPWR _21432_/X sky130_fd_sc_hd__or2_4
XFILLER_238_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15490__A1_N _14890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24151_ _24145_/CLK _18759_/Y HRESETn VGND VGND VPWR VPWR _24151_/Q sky130_fd_sc_hd__dfrtp_4
X_21363_ _13536_/A _12106_/A _12052_/Y _21580_/A VGND VGND VPWR VPWR _21363_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21852__B2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23102_ _24443_/Q _22851_/X _22108_/X _23101_/X VGND VGND VPWR VPWR _23102_/X sky130_fd_sc_hd__a211o_4
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20314_ _20314_/A VGND VGND VPWR VPWR _21666_/B sky130_fd_sc_hd__inv_2
X_24082_ _25365_/CLK _15497_/X HRESETn VGND VGND VPWR VPWR HREADYOUT sky130_fd_sc_hd__dfstp_4
X_21294_ _21122_/A VGND VGND VPWR VPWR _21295_/A sky130_fd_sc_hd__buf_2
XANTENNA__24583__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23033_ _16675_/Y _22842_/X _15592_/Y _22845_/X VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20245_ _18114_/B VGND VGND VPWR VPWR _20245_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20176_ _23490_/Q VGND VGND VPWR VPWR _20176_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16802__A1_N _16801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24984_ _24981_/CLK _15427_/X HRESETn VGND VGND VPWR VPWR _15162_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23935_ _24194_/CLK _23935_/D HRESETn VGND VGND VPWR VPWR _21002_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_217_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11880_ _17711_/B VGND VGND VPWR VPWR _11880_/Y sky130_fd_sc_hd__inv_2
X_23866_ _23628_/CLK _23866_/D VGND VGND VPWR VPWR _23866_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22828__A _22854_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22817_ _15012_/A _22673_/B _22816_/X VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23797_ _23445_/CLK _19298_/X VGND VGND VPWR VPWR _19297_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_199_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13550_ _13550_/A _17929_/A _24257_/Q VGND VGND VPWR VPWR _13550_/X sky130_fd_sc_hd__and3_4
XANTENNA__25300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22748_ _17341_/A _22437_/X _22747_/Y VGND VGND VPWR VPWR _22748_/X sky130_fd_sc_hd__o21a_4
X_25536_ _25539_/CLK _11828_/X HRESETn VGND VGND VPWR VPWR _11824_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_197_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21451__B _21450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16547__B1 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12501_ _12501_/A _12501_/B _12500_/Y VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__and3_4
XFILLER_241_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13481_ _13481_/A VGND VGND VPWR VPWR _13481_/X sky130_fd_sc_hd__buf_2
X_25467_ _25380_/CLK _12410_/X HRESETn VGND VGND VPWR VPWR _25467_/Q sky130_fd_sc_hd__dfrtp_4
X_22679_ _12439_/A _21542_/X _17762_/Y _22446_/A VGND VGND VPWR VPWR _22679_/X sky130_fd_sc_hd__o22a_4
XFILLER_157_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15220_ _15077_/D _15219_/X VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__or2_4
XANTENNA__13250__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12432_ _12424_/B VGND VGND VPWR VPWR _12432_/Y sky130_fd_sc_hd__inv_2
X_24418_ _24684_/CLK _16869_/X HRESETn VGND VGND VPWR VPWR _20102_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25398_ _24812_/CLK _25398_/D HRESETn VGND VGND VPWR VPWR _12899_/A sky130_fd_sc_hd__dfrtp_4
X_15151_ _25003_/Q VGND VGND VPWR VPWR _15345_/C sky130_fd_sc_hd__inv_2
X_12363_ _12363_/A VGND VGND VPWR VPWR _13038_/A sky130_fd_sc_hd__inv_2
X_24349_ _24354_/CLK _24349_/D HRESETn VGND VGND VPWR VPWR _17253_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_148_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21843__B2 _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14102_ _24014_/Q _14066_/A _14082_/X _14032_/A _14069_/B VGND VGND VPWR VPWR _14102_/X
+ sky130_fd_sc_hd__a32o_4
X_15082_ _15082_/A VGND VGND VPWR VPWR _15082_/Y sky130_fd_sc_hd__inv_2
X_12294_ _12294_/A _12247_/A _12293_/Y _12269_/Y VGND VGND VPWR VPWR _12296_/C sky130_fd_sc_hd__or4_4
XFILLER_154_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14033_ _14033_/A _14001_/X VGND VGND VPWR VPWR _14034_/D sky130_fd_sc_hd__or2_4
X_18910_ _23933_/Q VGND VGND VPWR VPWR _18910_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22399__A2 _22370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19890_ _19890_/A VGND VGND VPWR VPWR _21937_/B sky130_fd_sc_hd__inv_2
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ _16506_/A _24147_/Q _16506_/Y _18763_/A VGND VGND VPWR VPWR _18841_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15905__A _11830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18772_ _18772_/A _18772_/B VGND VGND VPWR VPWR _18773_/A sky130_fd_sc_hd__or2_4
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15984_ _12199_/Y _15983_/X _15905_/X _15983_/X VGND VGND VPWR VPWR _24763_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17723_ _24221_/Q VGND VGND VPWR VPWR _17723_/X sky130_fd_sc_hd__buf_2
X_14935_ _15076_/C VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__buf_2
XFILLER_76_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15038__B1 _25019_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17654_ _17641_/A _17651_/B _17653_/Y VGND VGND VPWR VPWR _24313_/D sky130_fd_sc_hd__and3_4
X_14866_ _14852_/X _14865_/Y _25052_/Q _14852_/X VGND VGND VPWR VPWR _14866_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16786__B1 _16530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16605_ _16603_/Y _16604_/X _16252_/X _16604_/X VGND VGND VPWR VPWR _24531_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21642__A _22387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13817_ _25276_/Q VGND VGND VPWR VPWR _13817_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22859__B1 _12350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12362__A2_N _24838_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17585_ _17701_/A _17529_/Y _17585_/C _17585_/D VGND VGND VPWR VPWR _17589_/B sky130_fd_sc_hd__or4_4
X_14797_ _18027_/A _14676_/X _18027_/A _14676_/X VGND VGND VPWR VPWR _14801_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19324_ _19323_/X VGND VGND VPWR VPWR _19324_/Y sky130_fd_sc_hd__inv_2
X_16536_ _24557_/Q VGND VGND VPWR VPWR _16536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ _13748_/A _14772_/A VGND VGND VPWR VPWR _13748_/X sky130_fd_sc_hd__or2_4
XANTENNA__16538__B1 _16537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19255_ _19253_/Y _19249_/X _19254_/X _19249_/A VGND VGND VPWR VPWR _19255_/X sky130_fd_sc_hd__a2bb2o_4
X_16467_ _15870_/B VGND VGND VPWR VPWR _16468_/A sky130_fd_sc_hd__buf_2
X_13679_ _23387_/Q _20834_/B VGND VGND VPWR VPWR _13679_/X sky130_fd_sc_hd__and2_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18206_ _18072_/X _18206_/B VGND VGND VPWR VPWR _18208_/B sky130_fd_sc_hd__or2_4
XFILLER_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15418_ _15398_/X VGND VGND VPWR VPWR _15419_/B sky130_fd_sc_hd__inv_2
X_19186_ _19186_/A VGND VGND VPWR VPWR _19186_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_23_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16398_ _16415_/A VGND VGND VPWR VPWR _16398_/X sky130_fd_sc_hd__buf_2
XANTENNA__20098__B1 _19761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18137_ _18169_/A _18135_/X _18136_/X VGND VGND VPWR VPWR _18137_/X sky130_fd_sc_hd__and3_4
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17567__A _24719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12575__B2 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15349_ _15303_/A _15352_/B _15348_/X VGND VGND VPWR VPWR _15349_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_145_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21089__A _15866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18068_ _18138_/A _18063_/X _18068_/C VGND VGND VPWR VPWR _18068_/X sky130_fd_sc_hd__or3_4
XFILLER_160_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16710__B1 _16613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17019_ _16028_/A _17057_/B _16033_/Y _24398_/Q VGND VGND VPWR VPWR _17020_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20030_ _20028_/Y _20029_/X _20007_/X _20029_/X VGND VGND VPWR VPWR _20030_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21817__A _21679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15277__B1 _15183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23339__B2 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_147_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _25316_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_239_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21981_ _23692_/Q _21981_/B _19605_/A _19608_/A VGND VGND VPWR VPWR _21981_/X sky130_fd_sc_hd__or4_4
XFILLER_227_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23720_ _23407_/CLK _23720_/D VGND VGND VPWR VPWR _23720_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ _20927_/X _20930_/X _16677_/A _20931_/X VGND VGND VPWR VPWR _20932_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16777__B1 _15759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _23644_/CLK _19723_/X VGND VGND VPWR VPWR _19722_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_214_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _20842_/A VGND VGND VPWR VPWR _20863_/X sky130_fd_sc_hd__buf_2
XFILLER_241_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22314__A2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22602_ _16519_/A _22440_/X _22545_/X VGND VGND VPWR VPWR _22602_/X sky130_fd_sc_hd__o21a_4
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _23582_/CLK _23582_/D VGND VGND VPWR VPWR _19919_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20794_ _20768_/B _20794_/B VGND VGND VPWR VPWR _20794_/Y sky130_fd_sc_hd__nor2_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25321_ _25316_/CLK _13508_/X HRESETn VGND VGND VPWR VPWR _12032_/A sky130_fd_sc_hd__dfrtp_4
X_22533_ _22533_/A _21604_/A VGND VGND VPWR VPWR _22534_/A sky130_fd_sc_hd__or2_4
XFILLER_210_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25252_ _25253_/CLK _13886_/X HRESETn VGND VGND VPWR VPWR _25252_/Q sky130_fd_sc_hd__dfrtp_4
X_22464_ _22459_/X _22461_/X _22462_/X _22463_/X VGND VGND VPWR VPWR _22464_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24764__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22383__A _22390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24203_ _24201_/CLK _18380_/X HRESETn VGND VGND VPWR VPWR _18376_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20089__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21415_ _14765_/X _20074_/Y VGND VGND VPWR VPWR _21415_/X sky130_fd_sc_hd__or2_4
X_25183_ _24112_/CLK _25183_/D HRESETn VGND VGND VPWR VPWR MSO_S2 sky130_fd_sc_hd__dfrtp_4
X_22395_ _22385_/A _19858_/Y _22209_/A VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__o21a_4
X_24134_ _24138_/CLK _24134_/D HRESETn VGND VGND VPWR VPWR _24134_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21346_ _24521_/Q _21341_/X _15676_/A _21345_/X VGND VGND VPWR VPWR _21347_/C sky130_fd_sc_hd__a211o_4
XFILLER_190_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13515__B1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24065_ _24500_/CLK _20917_/X HRESETn VGND VGND VPWR VPWR _20915_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19692__A _19048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21277_ _21277_/A _21269_/X _21277_/C VGND VGND VPWR VPWR _21277_/X sky130_fd_sc_hd__or3_4
XFILLER_104_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22830__B _22954_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23016_ _23016_/A VGND VGND VPWR VPWR _23016_/X sky130_fd_sc_hd__buf_2
X_20228_ _23470_/Q VGND VGND VPWR VPWR _21394_/B sky130_fd_sc_hd__inv_2
Xclkbuf_7_43_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_86_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20261__B1 _19769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20159_ _21924_/B _20156_/X _20112_/X _20156_/X VGND VGND VPWR VPWR _23497_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12981_ _12837_/Y _12984_/B _12875_/X VGND VGND VPWR VPWR _12981_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__25552__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24967_ _24966_/CLK _15466_/X HRESETn VGND VGND VPWR VPWR _13936_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_58_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22553__A2 _21320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14720_ _14719_/Y VGND VGND VPWR VPWR _22214_/A sky130_fd_sc_hd__buf_2
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13245__A _13320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _19626_/A VGND VGND VPWR VPWR _11932_/Y sky130_fd_sc_hd__inv_2
X_23918_ _23918_/CLK _23918_/D VGND VGND VPWR VPWR _23918_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_150_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24898_ _24651_/CLK _24898_/D HRESETn VGND VGND VPWR VPWR _15647_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11863_ _11859_/Y _11857_/X _11862_/X _11857_/X VGND VGND VPWR VPWR _25528_/D sky130_fd_sc_hd__a2bb2o_4
X_14651_ _18069_/A _14650_/X _18069_/A _14650_/X VGND VGND VPWR VPWR _14651_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23849_ _24100_/CLK _19155_/X VGND VGND VPWR VPWR _23849_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_233_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _17456_/A _11721_/A _11724_/A _13476_/D VGND VGND VPWR VPWR _13607_/B sky130_fd_sc_hd__or4_4
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17364_/A _17370_/B VGND VGND VPWR VPWR _17370_/X sky130_fd_sc_hd__or2_4
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11759_/X VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__buf_2
X_14582_ _14582_/A VGND VGND VPWR VPWR _14582_/Y sky130_fd_sc_hd__inv_2
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16321_ _16319_/Y _16320_/X _15963_/X _16320_/X VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ _13533_/A _13532_/X VGND VGND VPWR VPWR _13533_/X sky130_fd_sc_hd__and2_4
X_25519_ _25520_/CLK _25519_/D HRESETn VGND VGND VPWR VPWR _11887_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19040_ _19039_/Y _19037_/X _18969_/X _19037_/X VGND VGND VPWR VPWR _19040_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13464_ _13243_/X _13464_/B VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__or2_4
X_16252_ _16252_/A VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__buf_2
XFILLER_186_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23266__B1 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16940__B1 _16140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12415_ _12414_/X VGND VGND VPWR VPWR _12415_/Y sky130_fd_sc_hd__inv_2
X_15203_ _15203_/A _15202_/X VGND VGND VPWR VPWR _15203_/X sky130_fd_sc_hd__or2_4
XFILLER_173_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13395_ _13242_/X _13393_/X _13394_/X VGND VGND VPWR VPWR _13395_/X sky130_fd_sc_hd__and3_4
X_16183_ _14779_/A _14789_/A VGND VGND VPWR VPWR _16184_/B sky130_fd_sc_hd__and2_4
XANTENNA__20296__A2_N _20291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20525__B _20525_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23281__A3 _22291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17818__C _17562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12346_ _24843_/Q VGND VGND VPWR VPWR _12346_/Y sky130_fd_sc_hd__inv_2
X_15134_ _15134_/A VGND VGND VPWR VPWR _15134_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12309__B2 _24850_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15065_ _14893_/Y _14996_/X _15031_/X _15064_/X VGND VGND VPWR VPWR _15065_/X sky130_fd_sc_hd__o22a_4
X_19942_ _23573_/Q VGND VGND VPWR VPWR _19942_/Y sky130_fd_sc_hd__inv_2
X_12277_ _25466_/Q _12264_/Y _12263_/Y _24757_/Q VGND VGND VPWR VPWR _12280_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12324__A _24844_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14016_ _25244_/Q VGND VGND VPWR VPWR _14021_/B sky130_fd_sc_hd__buf_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22241__A1 _13560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19873_ _19873_/A VGND VGND VPWR VPWR _19873_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20252__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18824_ _18689_/B _18824_/B VGND VGND VPWR VPWR _18824_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15635__A _15626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18011__A _18098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18755_ _24152_/Q _18755_/B VGND VGND VPWR VPWR _18757_/B sky130_fd_sc_hd__or2_4
XANTENNA__25293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_0_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_15967_ HWDATA[19] VGND VGND VPWR VPWR _15967_/X sky130_fd_sc_hd__buf_2
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14482__B2 _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _24297_/Q _17705_/Y VGND VGND VPWR VPWR _17706_/X sky130_fd_sc_hd__or2_4
XFILLER_208_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13155__A _13212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14918_ _15256_/A _24419_/Q _15256_/A _24419_/Q VGND VGND VPWR VPWR _14918_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18686_ _18686_/A VGND VGND VPWR VPWR _18687_/D sky130_fd_sc_hd__inv_2
XFILLER_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16759__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15898_ _15894_/X _15895_/X _16238_/A _22755_/A _15896_/X VGND VGND VPWR VPWR _24805_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17637_ _17579_/B _17636_/X VGND VGND VPWR VPWR _17637_/X sky130_fd_sc_hd__or2_4
X_14849_ _24005_/D _14848_/Y _25202_/Q _24005_/D VGND VGND VPWR VPWR _25057_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21091__B _21091_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17568_ _17567_/Y VGND VGND VPWR VPWR _17663_/A sky130_fd_sc_hd__buf_2
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15982__A1 _15797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19307_ _23794_/Q VGND VGND VPWR VPWR _19307_/Y sky130_fd_sc_hd__inv_2
X_16519_ _16519_/A VGND VGND VPWR VPWR _16519_/Y sky130_fd_sc_hd__inv_2
X_17499_ _17470_/X _17480_/X _17499_/C _17498_/X VGND VGND VPWR VPWR _17499_/X sky130_fd_sc_hd__or4_4
X_19238_ _13220_/B VGND VGND VPWR VPWR _19238_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20716__A _20716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19169_ _19032_/A VGND VGND VPWR VPWR _19169_/X sky130_fd_sc_hd__buf_2
XFILLER_192_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21200_ _21182_/A _21200_/B VGND VGND VPWR VPWR _21200_/X sky130_fd_sc_hd__or2_4
XFILLER_145_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22180_ _22179_/Y _21353_/X _14137_/Y _14229_/A VGND VGND VPWR VPWR _22181_/A sky130_fd_sc_hd__o22a_4
XFILLER_219_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22931__A _22694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21131_ _21047_/X _21128_/X _21129_/X _21130_/Y VGND VGND VPWR VPWR _21132_/C sky130_fd_sc_hd__a211o_4
X_21062_ _21062_/A VGND VGND VPWR VPWR _21063_/A sky130_fd_sc_hd__buf_2
XANTENNA__21547__A _21126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20013_ _21187_/B _20006_/X _19900_/X _19988_/Y VGND VGND VPWR VPWR _23549_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24821_ _24856_/CLK _24821_/D HRESETn VGND VGND VPWR VPWR _24821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21964_ _21949_/A _21962_/X _21964_/C VGND VGND VPWR VPWR _21964_/X sky130_fd_sc_hd__and3_4
X_24752_ _24735_/CLK _16007_/X HRESETn VGND VGND VPWR VPWR _15999_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_242_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20915_ _24064_/Q _20915_/B _24063_/Q _20907_/B VGND VGND VPWR VPWR _20915_/X sky130_fd_sc_hd__or4_4
X_23703_ _23703_/CLK _19567_/X VGND VGND VPWR VPWR _19564_/A sky130_fd_sc_hd__dfxtp_4
X_24683_ _24657_/CLK _16198_/X HRESETn VGND VGND VPWR VPWR _23341_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_161_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _21267_/A VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__buf_2
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _23644_/CLK _23634_/D VGND VGND VPWR VPWR _13299_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _24050_/Q VGND VGND VPWR VPWR _20846_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16095__B _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19164__B2 _19159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _23565_/CLK _19963_/X VGND VGND VPWR VPWR _19962_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_168_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20777_ _20775_/Y _20772_/X _20776_/X VGND VGND VPWR VPWR _20777_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22516_ _21596_/A _22516_/B VGND VGND VPWR VPWR _22516_/Y sky130_fd_sc_hd__nor2_4
X_25304_ _24913_/CLK _13681_/X HRESETn VGND VGND VPWR VPWR _25304_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_210_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23496_ _23513_/CLK _23496_/D VGND VGND VPWR VPWR _23496_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__B2 _24860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22447_ _22447_/A VGND VGND VPWR VPWR _22732_/A sky130_fd_sc_hd__buf_2
X_25235_ _25246_/CLK _25235_/D HRESETn VGND VGND VPWR VPWR _13992_/A sky130_fd_sc_hd__dfrtp_4
X_12200_ _12200_/A VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__inv_2
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13180_ _13199_/A _23620_/Q VGND VGND VPWR VPWR _13181_/C sky130_fd_sc_hd__or2_4
X_25166_ _24121_/CLK _14367_/X HRESETn VGND VGND VPWR VPWR MSO_S3 sky130_fd_sc_hd__dfrtp_4
XANTENNA__22471__A1 _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22378_ _22085_/A _19277_/Y VGND VGND VPWR VPWR _22380_/B sky130_fd_sc_hd__or2_4
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22471__B2 _22470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12131_ _12175_/A _12128_/X _11871_/X _12128_/X VGND VGND VPWR VPWR _25475_/D sky130_fd_sc_hd__a2bb2o_4
X_24117_ _25145_/CLK _24117_/D HRESETn VGND VGND VPWR VPWR _24117_/Q sky130_fd_sc_hd__dfrtp_4
X_21329_ _15134_/A _22945_/A VGND VGND VPWR VPWR _21338_/B sky130_fd_sc_hd__or2_4
XFILLER_163_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25097_ _25093_/CLK _14602_/X HRESETn VGND VGND VPWR VPWR _25097_/Q sky130_fd_sc_hd__dfrtp_4
X_12062_ _16378_/A _11721_/Y _16190_/C _13476_/D VGND VGND VPWR VPWR _21583_/B sky130_fd_sc_hd__or4_4
X_24048_ _24485_/CLK _24048_/D HRESETn VGND VGND VPWR VPWR _24048_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21457__A _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16870_ _20105_/A VGND VGND VPWR VPWR _16870_/X sky130_fd_sc_hd__buf_2
XFILLER_150_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15149__A2_N _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15821_ _15818_/A VGND VGND VPWR VPWR _15821_/X sky130_fd_sc_hd__buf_2
XFILLER_93_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15174__B _15294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_130_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23735_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18540_ _18540_/A _18540_/B _18543_/A _18543_/B VGND VGND VPWR VPWR _18540_/X sky130_fd_sc_hd__or4_4
X_15752_ HWDATA[15] VGND VGND VPWR VPWR _15752_/X sky130_fd_sc_hd__buf_2
XFILLER_206_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12964_ _12855_/A _12961_/X VGND VGND VPWR VPWR _12964_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_193_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24485_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_205_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14703_ _18914_/A _13759_/Y _13767_/B VGND VGND VPWR VPWR _14703_/X sky130_fd_sc_hd__a21o_4
XFILLER_218_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11915_ _11881_/X _11914_/X _11905_/X _11913_/A VGND VGND VPWR VPWR _25521_/D sky130_fd_sc_hd__a22oi_4
X_18471_ _18471_/A _18543_/A _18539_/A _18471_/D VGND VGND VPWR VPWR _18472_/C sky130_fd_sc_hd__or4_4
XFILLER_205_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15683_ _16382_/A VGND VGND VPWR VPWR _15683_/X sky130_fd_sc_hd__buf_2
X_12895_ _12825_/Y _12895_/B _12609_/X VGND VGND VPWR VPWR _12895_/X sky130_fd_sc_hd__or3_4
X_17422_ _17422_/A VGND VGND VPWR VPWR _21373_/A sky130_fd_sc_hd__buf_2
XFILLER_233_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14634_ _14633_/X VGND VGND VPWR VPWR _14634_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11846_ HWDATA[6] VGND VGND VPWR VPWR _11847_/A sky130_fd_sc_hd__buf_2
XFILLER_233_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24686__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17353_/A VGND VGND VPWR VPWR _17363_/A sky130_fd_sc_hd__buf_2
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11759_/X VGND VGND VPWR VPWR _11777_/X sky130_fd_sc_hd__buf_2
X_14565_ _14564_/X VGND VGND VPWR VPWR _14595_/A sky130_fd_sc_hd__inv_2
XFILLER_186_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24615__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _24643_/Q VGND VGND VPWR VPWR _16304_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13516_ _13516_/A VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__buf_2
X_17284_ _17286_/B VGND VGND VPWR VPWR _17284_/Y sky130_fd_sc_hd__inv_2
X_14496_ _25121_/Q VGND VGND VPWR VPWR _14496_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19023_ _19022_/Y _19020_/X _18908_/X _19020_/X VGND VGND VPWR VPWR _19023_/X sky130_fd_sc_hd__a2bb2o_4
X_16235_ _16264_/A VGND VGND VPWR VPWR _16235_/X sky130_fd_sc_hd__buf_2
X_13447_ _13310_/X _13445_/X _13446_/X VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__and3_4
XFILLER_173_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18006__A _18006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13378_ _13410_/A _23871_/Q VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__or2_4
X_16166_ _16166_/A VGND VGND VPWR VPWR _16166_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ _25010_/Q VGND VGND VPWR VPWR _15318_/C sky130_fd_sc_hd__inv_2
X_12329_ _12329_/A VGND VGND VPWR VPWR _12329_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16097_ _16096_/X VGND VGND VPWR VPWR _16097_/X sky130_fd_sc_hd__buf_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14152__B1 _25145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15048_ _15248_/A _16776_/A _15248_/A _16776_/A VGND VGND VPWR VPWR _15049_/D sky130_fd_sc_hd__a2bb2o_4
X_19925_ _19925_/A VGND VGND VPWR VPWR _19925_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14988__A2_N _14976_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19856_ _20146_/A VGND VGND VPWR VPWR _19856_/X sky130_fd_sc_hd__buf_2
XANTENNA__25403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18807_ _18799_/B _18799_/C _18729_/X _18803_/Y VGND VGND VPWR VPWR _18808_/A sky130_fd_sc_hd__a211o_4
X_19787_ _19837_/A _13771_/X _19278_/X VGND VGND VPWR VPWR _19788_/A sky130_fd_sc_hd__or3_4
X_16999_ _16972_/X _16980_/X _16989_/X _16998_/X VGND VGND VPWR VPWR _17027_/A sky130_fd_sc_hd__or4_4
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19918__B1 _19643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18738_ _18681_/Y _18736_/A VGND VGND VPWR VPWR _18739_/C sky130_fd_sc_hd__or2_4
XFILLER_209_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18669_ _16556_/Y _24161_/Q _16556_/Y _24161_/Q VGND VGND VPWR VPWR _18673_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20700_ _20699_/X VGND VGND VPWR VPWR _20700_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21680_ _17738_/A VGND VGND VPWR VPWR _22274_/A sky130_fd_sc_hd__buf_2
XFILLER_240_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22926__A _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20631_ _20631_/A VGND VGND VPWR VPWR _23988_/D sky130_fd_sc_hd__inv_2
XANTENNA__21830__A _21815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17223__A2_N _17212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23350_ _23331_/X _23334_/X _23338_/Y _23349_/X VGND VGND VPWR VPWR HRDATA[31] sky130_fd_sc_hd__a211o_4
X_20562_ _14453_/Y _20551_/X _20608_/A _20561_/X VGND VGND VPWR VPWR _20563_/A sky130_fd_sc_hd__a211o_4
XFILLER_149_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22301_ _21604_/A _22301_/B VGND VGND VPWR VPWR _22301_/Y sky130_fd_sc_hd__nor2_4
XFILLER_164_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23281_ _12791_/Y _22725_/X _22291_/B _12555_/Y _22862_/X VGND VGND VPWR VPWR _23281_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_192_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20493_ _23978_/Q _24093_/Q VGND VGND VPWR VPWR _20493_/X sky130_fd_sc_hd__and2_4
XFILLER_20_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25020_ _25018_/CLK _15278_/X HRESETn VGND VGND VPWR VPWR _25020_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22232_ _21260_/A _22230_/X _22231_/X VGND VGND VPWR VPWR _22236_/B sky130_fd_sc_hd__and3_4
XFILLER_118_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22661__A _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22163_ _22146_/B _22162_/X _22986_/A _25530_/Q _22947_/A VGND VGND VPWR VPWR _22163_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_246_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21114_ _16000_/X VGND VGND VPWR VPWR _21321_/A sky130_fd_sc_hd__buf_2
XANTENNA__14143__B1 _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18409__B1 _23218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22094_ _22094_/A _22094_/B VGND VGND VPWR VPWR _22094_/X sky130_fd_sc_hd__or2_4
XANTENNA__12899__A _12899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15891__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21045_ _21045_/A _14484_/A VGND VGND VPWR VPWR _21046_/A sky130_fd_sc_hd__or2_4
XFILLER_115_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24804_ _24794_/CLK _15899_/X HRESETn VGND VGND VPWR VPWR _22726_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17490__A _24328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_203_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _23973_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21716__B1 _24828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22996_ _22787_/X _22992_/Y _22881_/X _22995_/X VGND VGND VPWR VPWR _22996_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_215_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24735_ _24735_/CLK _16050_/X HRESETn VGND VGND VPWR VPWR _24735_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_9_0_HCLK clkbuf_8_9_0_HCLK/A VGND VGND VPWR VPWR _23684_/CLK sky130_fd_sc_hd__clkbuf_1
X_21947_ _21947_/A _19974_/Y VGND VGND VPWR VPWR _21949_/B sky130_fd_sc_hd__or2_4
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11700_/A VGND VGND VPWR VPWR _13698_/A sky130_fd_sc_hd__inv_2
XFILLER_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A _12680_/B _12680_/C VGND VGND VPWR VPWR _12680_/X sky130_fd_sc_hd__and3_4
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _24423_/Q _22299_/B _21741_/A _21877_/X VGND VGND VPWR VPWR _21878_/X sky130_fd_sc_hd__a211o_4
X_24666_ _24666_/CLK _16243_/X HRESETn VGND VGND VPWR VPWR _22716_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22836__A _22836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _23386_/D _13147_/A _13147_/B _23336_/A _20744_/A VGND VGND VPWR VPWR _20829_/X
+ sky130_fd_sc_hd__a32o_4
X_23617_ _25507_/CLK _19825_/X VGND VGND VPWR VPWR _23617_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24597_ _24601_/CLK _24597_/D HRESETn VGND VGND VPWR VPWR _16432_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14350_ _14350_/A VGND VGND VPWR VPWR _14350_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22692__A1 _21113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23548_ _23563_/CLK _23548_/D VGND VGND VPWR VPWR _23548_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13177_/A _13299_/X _13301_/C VGND VGND VPWR VPWR _13301_/X sky130_fd_sc_hd__and3_4
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _14279_/Y _14280_/X _13812_/X _14280_/X VGND VGND VPWR VPWR _25192_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23479_ _23494_/CLK _23479_/D VGND VGND VPWR VPWR _20204_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ _13387_/A _13229_/X _13231_/X VGND VGND VPWR VPWR _13239_/B sky130_fd_sc_hd__and3_4
X_16020_ _16018_/Y _16019_/X _11770_/X _16019_/X VGND VGND VPWR VPWR _24747_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25218_ _25215_/CLK _25218_/D HRESETn VGND VGND VPWR VPWR _14107_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__22571__A _16348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13163_ _13177_/A _13158_/X _13162_/X VGND VGND VPWR VPWR _13163_/X sky130_fd_sc_hd__and3_4
X_25149_ _25223_/CLK _14424_/X HRESETn VGND VGND VPWR VPWR _25149_/Q sky130_fd_sc_hd__dfstp_4
X_12114_ _12113_/Y _12111_/X _11838_/X _12111_/X VGND VGND VPWR VPWR _25482_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13094_ _12326_/Y _13106_/B VGND VGND VPWR VPWR _13104_/B sky130_fd_sc_hd__or2_4
X_17971_ _17973_/A VGND VGND VPWR VPWR _18031_/A sky130_fd_sc_hd__inv_2
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19710_ _19710_/A VGND VGND VPWR VPWR _19710_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22747__A2 _21320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15882__B1 _23162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12045_ _25497_/Q VGND VGND VPWR VPWR _12045_/Y sky130_fd_sc_hd__inv_2
X_16922_ _16922_/A _16922_/B _16922_/C _16921_/X VGND VGND VPWR VPWR _16922_/X sky130_fd_sc_hd__or4_4
XANTENNA__19073__B1 _18999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19641_ _19641_/A VGND VGND VPWR VPWR _21695_/B sky130_fd_sc_hd__inv_2
XFILLER_238_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16853_ _16853_/A VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__buf_2
XFILLER_120_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23157__C1 _23156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15804_ _15796_/X VGND VGND VPWR VPWR _15804_/X sky130_fd_sc_hd__buf_2
XFILLER_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19572_ _23700_/Q VGND VGND VPWR VPWR _22360_/B sky130_fd_sc_hd__inv_2
X_16784_ _15017_/Y _16782_/X _16613_/X _16782_/X VGND VGND VPWR VPWR _16784_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13996_ _25247_/Q VGND VGND VPWR VPWR _14062_/A sky130_fd_sc_hd__buf_2
XANTENNA__24867__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18523_ _24186_/Q _18523_/B VGND VGND VPWR VPWR _18524_/C sky130_fd_sc_hd__or2_4
X_15735_ _15557_/X _15722_/X _15734_/X _24885_/Q _15720_/X VGND VGND VPWR VPWR _15735_/X
+ sky130_fd_sc_hd__a32o_4
X_12947_ _12947_/A VGND VGND VPWR VPWR _12947_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17387__B1 _17280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18454_ _23250_/A _18445_/Y _16268_/Y _24167_/Q VGND VGND VPWR VPWR _18456_/C sky130_fd_sc_hd__a2bb2o_4
X_15666_ _21105_/B VGND VGND VPWR VPWR _15667_/A sky130_fd_sc_hd__buf_2
XANTENNA__15937__A1 _15678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12878_ _12878_/A _12865_/X VGND VGND VPWR VPWR _12878_/X sky130_fd_sc_hd__or2_4
XFILLER_222_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17405_/A _20661_/A VGND VGND VPWR VPWR _17406_/B sky130_fd_sc_hd__or2_4
X_14617_ _13575_/Y _14570_/B VGND VGND VPWR VPWR _14617_/Y sky130_fd_sc_hd__nand2_4
X_11829_ _25535_/Q VGND VGND VPWR VPWR _11829_/Y sky130_fd_sc_hd__inv_2
X_18385_ _18383_/Y _18379_/X _18386_/A _18384_/X VGND VGND VPWR VPWR _24201_/D sky130_fd_sc_hd__a2bb2o_4
X_15597_ _15614_/A VGND VGND VPWR VPWR _15597_/X sky130_fd_sc_hd__buf_2
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17336_ _17262_/Y _17326_/D _17288_/X _17333_/Y VGND VGND VPWR VPWR _17336_/X sky130_fd_sc_hd__a211o_4
X_14548_ _14548_/A VGND VGND VPWR VPWR _14548_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11888__A _11889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17267_ _17245_/Y _17267_/B VGND VGND VPWR VPWR _17267_/X sky130_fd_sc_hd__or2_4
X_14479_ _14479_/A VGND VGND VPWR VPWR _14479_/X sky130_fd_sc_hd__buf_2
XANTENNA__14264__A _14264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19006_ _23899_/Q VGND VGND VPWR VPWR _19006_/Y sky130_fd_sc_hd__inv_2
X_16218_ _16217_/Y _16215_/X _11780_/X _16215_/X VGND VGND VPWR VPWR _16218_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18639__B1 _16608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17198_ _17197_/Y VGND VGND VPWR VPWR _17198_/X sky130_fd_sc_hd__buf_2
X_16149_ _16147_/Y _16148_/X _11827_/X _16148_/X VGND VGND VPWR VPWR _24697_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19908_ _22255_/B _19905_/X _19629_/X _19905_/X VGND VGND VPWR VPWR _23587_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13608__A _14679_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19064__B1 _18969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21825__A _21687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18811__B1 _18714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19839_ _19838_/Y VGND VGND VPWR VPWR _19839_/X sky130_fd_sc_hd__buf_2
XFILLER_229_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22850_ _24602_/Q _22849_/X VGND VGND VPWR VPWR _22856_/B sky130_fd_sc_hd__or2_4
XANTENNA__21544__B _22897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21801_ _21800_/X VGND VGND VPWR VPWR _21801_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22781_ _22487_/A _22780_/X VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__and2_4
XANTENNA__21174__A1 _16801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14439__A _25143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21732_ _14277_/Y _21375_/X VGND VGND VPWR VPWR _21732_/Y sky130_fd_sc_hd__nor2_4
X_24520_ _24552_/CLK _16632_/X HRESETn VGND VGND VPWR VPWR _16631_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_33_0_HCLK clkbuf_8_33_0_HCLK/A VGND VGND VPWR VPWR _23488_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20921__A1 _16682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16050__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_96_0_HCLK clkbuf_8_97_0_HCLK/A VGND VGND VPWR VPWR _24726_/CLK sky130_fd_sc_hd__clkbuf_1
X_21663_ _21662_/X VGND VGND VPWR VPWR _21663_/Y sky130_fd_sc_hd__inv_2
X_24451_ _25011_/CLK _16802_/X HRESETn VGND VGND VPWR VPWR _24451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_212_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22123__B1 _21064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20614_ _20614_/A _20609_/B VGND VGND VPWR VPWR _20614_/X sky130_fd_sc_hd__or2_4
X_23402_ _23400_/CLK _23402_/D VGND VGND VPWR VPWR _23402_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24382_ _24407_/CLK _17162_/Y HRESETn VGND VGND VPWR VPWR _17051_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22674__A1 _15718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21594_ _16627_/Y _21588_/X _21591_/X _21593_/X VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22674__B2 _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23333_ _17274_/A _22493_/X _25404_/Q _22453_/X VGND VGND VPWR VPWR _23333_/X sky130_fd_sc_hd__a2bb2o_4
X_20545_ _20446_/C _20513_/X _20461_/D _14504_/X _20451_/X VGND VGND VPWR VPWR _20545_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_119_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17550__B1 _25553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23264_ _24375_/Q _21034_/X VGND VGND VPWR VPWR _23267_/B sky130_fd_sc_hd__or2_4
X_20476_ _20455_/B _20476_/B _20476_/C _20476_/D VGND VGND VPWR VPWR _20476_/X sky130_fd_sc_hd__or4_4
XANTENNA__25396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22215_ _22210_/A _20174_/Y VGND VGND VPWR VPWR _22217_/B sky130_fd_sc_hd__or2_4
X_25003_ _25002_/CLK _25003_/D HRESETn VGND VGND VPWR VPWR _25003_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23195_ _23173_/X _23176_/X _23180_/Y _23194_/X VGND VGND VPWR VPWR HRDATA[26] sky130_fd_sc_hd__a211o_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21719__B _21719_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22146_ _15634_/A _22146_/B VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__or2_4
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22077_ _22392_/A _22077_/B VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__or2_4
XANTENNA__17066__C1 _17065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21028_ _21027_/X VGND VGND VPWR VPWR _21029_/A sky130_fd_sc_hd__inv_2
XFILLER_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13850_ _13552_/Y _13848_/X _13849_/X _13848_/X VGND VGND VPWR VPWR _13850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _24807_/Q VGND VGND VPWR VPWR _12801_/Y sky130_fd_sc_hd__inv_2
X_13781_ _13781_/A VGND VGND VPWR VPWR _16464_/A sky130_fd_sc_hd__buf_2
XANTENNA__21173__C _21173_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21165__A1 _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _22956_/X _22979_/B _22979_/C _22978_/X VGND VGND VPWR VPWR HRDATA[20] sky130_fd_sc_hd__or4_4
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15520_ _15503_/A VGND VGND VPWR VPWR _15520_/X sky130_fd_sc_hd__buf_2
XANTENNA__18030__A1 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12732_ _12732_/A VGND VGND VPWR VPWR _12733_/B sky130_fd_sc_hd__inv_2
X_24718_ _24651_/CLK _24718_/D HRESETn VGND VGND VPWR VPWR _24718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16041__B1 _15972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21470__A _21815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15451_ _14289_/X _24085_/Q _15450_/Y _13942_/X _15447_/X VGND VGND VPWR VPWR _15451_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_230_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12663_ _12616_/A _12666_/B _12662_/X VGND VGND VPWR VPWR _12663_/Y sky130_fd_sc_hd__a21oi_4
X_24649_ _24015_/CLK _16286_/X HRESETn VGND VGND VPWR VPWR _24649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22285__B _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _25154_/Q VGND VGND VPWR VPWR _14402_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18138_/A _18170_/B _18170_/C VGND VGND VPWR VPWR _18171_/C sky130_fd_sc_hd__or3_4
Xclkbuf_5_4_0_HCLK clkbuf_5_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15369_/X VGND VGND VPWR VPWR _15383_/B sky130_fd_sc_hd__inv_2
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12630_/A _24886_/Q _25426_/Q _12593_/Y VGND VGND VPWR VPWR _12594_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _17106_/A _17115_/B _17120_/Y VGND VGND VPWR VPWR _24394_/D sky130_fd_sc_hd__and3_4
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _14338_/A _25175_/Q _25174_/Q VGND VGND VPWR VPWR _25175_/D sky130_fd_sc_hd__a21o_4
XFILLER_183_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17541__B1 _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _24378_/Q VGND VGND VPWR VPWR _17052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22417__A1 _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14264_ _14264_/A VGND VGND VPWR VPWR _21375_/A sky130_fd_sc_hd__buf_2
XANTENNA__22417__B2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16003_ _16003_/A _16288_/B VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__and2_4
XANTENNA__20428__B1 _11851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13215_ _13450_/A _13215_/B VGND VGND VPWR VPWR _13216_/C sky130_fd_sc_hd__or2_4
XANTENNA__25066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ _14194_/Y VGND VGND VPWR VPWR _20504_/A sky130_fd_sc_hd__buf_2
XFILLER_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13146_ _20822_/A _20822_/B _24045_/Q _13145_/X VGND VGND VPWR VPWR _13147_/B sky130_fd_sc_hd__or4_4
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15855__B1 _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13077_ _12997_/D _13061_/B _13019_/A _13074_/Y VGND VGND VPWR VPWR _13077_/X sky130_fd_sc_hd__a211o_4
X_17954_ _17954_/A _17954_/B _17954_/C VGND VGND VPWR VPWR _17954_/X sky130_fd_sc_hd__or3_4
X_12028_ _24109_/Q _12024_/X VGND VGND VPWR VPWR _12030_/A sky130_fd_sc_hd__and2_4
X_16905_ _16134_/Y _17767_/A _16134_/Y _17767_/A VGND VGND VPWR VPWR _16913_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17885_ _17757_/C _17858_/X _17798_/X _17883_/B VGND VGND VPWR VPWR _17886_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16739__A _16738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15607__B1 _11805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16836_ _24434_/Q VGND VGND VPWR VPWR _16836_/Y sky130_fd_sc_hd__inv_2
X_19624_ _19623_/X VGND VGND VPWR VPWR _19624_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15083__B2 _16434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19555_ _19554_/Y _19552_/X _19418_/X _19552_/X VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__a2bb2o_4
X_16767_ _16737_/Y VGND VGND VPWR VPWR _16782_/A sky130_fd_sc_hd__buf_2
X_13979_ _13949_/Y _13953_/Y _13978_/X _13979_/D VGND VGND VPWR VPWR _13980_/A sky130_fd_sc_hd__or4_4
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24630__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18506_ _18445_/Y _18504_/X _18505_/X _18500_/B VGND VGND VPWR VPWR _18507_/A sky130_fd_sc_hd__a211o_4
X_15718_ _15718_/A _15854_/B VGND VGND VPWR VPWR _15725_/A sky130_fd_sc_hd__or2_4
XFILLER_179_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19486_ _23731_/Q VGND VGND VPWR VPWR _22244_/B sky130_fd_sc_hd__inv_2
X_16698_ _16696_/Y _16692_/X _15756_/X _16697_/X VGND VGND VPWR VPWR _16698_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12841__B1 _12828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16032__B1 _15963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22476__A _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18437_ _16240_/Y _24177_/Q _16240_/Y _24177_/Q VGND VGND VPWR VPWR _18438_/D sky130_fd_sc_hd__a2bb2o_4
X_15649_ _17456_/A _11721_/Y _16190_/C _15559_/D VGND VGND VPWR VPWR _22121_/A sky130_fd_sc_hd__or4_4
XANTENNA__22907__C _22900_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18368_ _18368_/A VGND VGND VPWR VPWR _18368_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21459__A2 _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17319_ _17229_/Y _17318_/X VGND VGND VPWR VPWR _17322_/B sky130_fd_sc_hd__or2_4
XFILLER_147_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18299_ _21210_/A VGND VGND VPWR VPWR _18300_/B sky130_fd_sc_hd__buf_2
XFILLER_135_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20330_ _20328_/Y _20324_/X _19996_/X _20329_/X VGND VGND VPWR VPWR _23433_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22959__A2 _21039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _20260_/Y _20258_/X _19769_/X _20258_/X VGND VGND VPWR VPWR _23459_/D sky130_fd_sc_hd__a2bb2o_4
X_22000_ _21520_/X _21929_/X _21969_/X _21984_/Y _21999_/Y VGND VGND VPWR VPWR _22000_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16099__B1 _11752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20192_ _20191_/X VGND VGND VPWR VPWR _20193_/A sky130_fd_sc_hd__inv_2
XFILLER_143_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15846__B1 _24828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24340__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24789__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23951_ _23960_/CLK _23951_/D HRESETn VGND VGND VPWR VPWR _23951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_243_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24718__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16649__A _15565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19849__A2_N _19844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22902_ _24603_/Q _15681_/X VGND VGND VPWR VPWR _22906_/B sky130_fd_sc_hd__or2_4
XFILLER_96_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15553__A _22575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23882_ _23880_/CLK _23882_/D VGND VGND VPWR VPWR _19060_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_217_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22833_ _17212_/A _21065_/X VGND VGND VPWR VPWR _22836_/B sky130_fd_sc_hd__or2_4
XFILLER_244_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25552_ _24697_/CLK _11767_/X HRESETn VGND VGND VPWR VPWR _25552_/Q sky130_fd_sc_hd__dfrtp_4
X_22764_ _22562_/X _22763_/X _22157_/C _25540_/Q _22940_/A VGND VGND VPWR VPWR _22764_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22386__A _22090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _24503_/CLK _24503_/D HRESETn VGND VGND VPWR VPWR _16682_/A sky130_fd_sc_hd__dfrtp_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21715_ _21715_/A _22897_/A VGND VGND VPWR VPWR _21715_/X sky130_fd_sc_hd__or2_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22695_ _16696_/Y _22695_/B VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__and2_4
X_25483_ _25316_/CLK _25483_/D HRESETn VGND VGND VPWR VPWR _25483_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16384__A _16384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21646_ _21646_/A _21644_/X _21646_/C VGND VGND VPWR VPWR _21646_/X sky130_fd_sc_hd__and3_4
X_24434_ _24431_/CLK _24434_/D HRESETn VGND VGND VPWR VPWR _24434_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21577_ _21577_/A _21577_/B VGND VGND VPWR VPWR _21577_/X sky130_fd_sc_hd__or2_4
X_24365_ _24346_/CLK _17328_/X HRESETn VGND VGND VPWR VPWR _24365_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22833__B _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20528_ _20448_/X _20461_/D VGND VGND VPWR VPWR _20528_/X sky130_fd_sc_hd__and2_4
X_23316_ _23188_/X _23313_/X _23315_/X VGND VGND VPWR VPWR _23317_/D sky130_fd_sc_hd__and3_4
XFILLER_165_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24296_ _25528_/CLK _17709_/Y HRESETn VGND VGND VPWR VPWR _24296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23010__A _24673_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20459_ _25116_/Q _14510_/B _25117_/Q VGND VGND VPWR VPWR _20460_/A sky130_fd_sc_hd__or3_4
X_23247_ _23136_/X _23247_/B VGND VGND VPWR VPWR _23247_/Y sky130_fd_sc_hd__nor2_4
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13000_ _12339_/Y _12326_/Y _12332_/Y _12386_/Y VGND VGND VPWR VPWR _13005_/A sky130_fd_sc_hd__or4_4
XFILLER_134_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17826__A1 _16950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23178_ _15581_/Y _23140_/B VGND VGND VPWR VPWR _23178_/X sky130_fd_sc_hd__and2_4
XFILLER_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21168__C _21173_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15837__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22129_ _22129_/A _22129_/B VGND VGND VPWR VPWR _22129_/X sky130_fd_sc_hd__and2_4
XANTENNA__21465__A _21210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14951_ _15282_/A VGND VGND VPWR VPWR _15275_/A sky130_fd_sc_hd__inv_2
XFILLER_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13902_ _13902_/A _13924_/C _13944_/A _15435_/B VGND VGND VPWR VPWR _13902_/X sky130_fd_sc_hd__or4_4
XFILLER_236_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17670_ _17670_/A VGND VGND VPWR VPWR _24308_/D sky130_fd_sc_hd__inv_2
XANTENNA__24125__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14882_ _14878_/Y _14881_/Y _14873_/X VGND VGND VPWR VPWR _14882_/X sky130_fd_sc_hd__o21a_4
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16262__B1 _16066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16621_ _16620_/Y _16618_/X _16537_/X _16618_/X VGND VGND VPWR VPWR _24525_/D sky130_fd_sc_hd__a2bb2o_4
X_13833_ _13571_/Y _13831_/X _11813_/X _13831_/X VGND VGND VPWR VPWR _13833_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19340_ _18177_/B VGND VGND VPWR VPWR _19340_/Y sky130_fd_sc_hd__inv_2
X_16552_ _16552_/A _16468_/B VGND VGND VPWR VPWR _16623_/A sky130_fd_sc_hd__nor2_4
X_13764_ _18914_/A _13761_/X _13762_/X _14706_/A VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__or4_4
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12823__B1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22296__A _21606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15503_ _15503_/A VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__buf_2
X_12715_ _12550_/Y _12731_/A VGND VGND VPWR VPWR _12715_/X sky130_fd_sc_hd__or2_4
X_19271_ _19258_/Y VGND VGND VPWR VPWR _19271_/X sky130_fd_sc_hd__buf_2
X_16483_ _16495_/A VGND VGND VPWR VPWR _16483_/X sky130_fd_sc_hd__buf_2
X_13695_ _11672_/Y _13695_/B VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__or2_4
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16294__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18222_ _18158_/A _19072_/A VGND VGND VPWR VPWR _18222_/X sky130_fd_sc_hd__or2_4
X_15434_ _15433_/X VGND VGND VPWR VPWR _15434_/Y sky130_fd_sc_hd__inv_2
X_12646_ _12636_/A _12646_/B _12645_/X VGND VGND VPWR VPWR _12646_/X sky130_fd_sc_hd__and3_4
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _18084_/X _18994_/A VGND VGND VPWR VPWR _18154_/C sky130_fd_sc_hd__or2_4
X_15365_ _15365_/A _15363_/A VGND VGND VPWR VPWR _15366_/C sky130_fd_sc_hd__or2_4
XANTENNA__25247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12577_ _12618_/D _24874_/Q _12618_/D _24874_/Q VGND VGND VPWR VPWR _12577_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17104_ _24399_/Q _17104_/B VGND VGND VPWR VPWR _17104_/X sky130_fd_sc_hd__or2_4
X_14316_ _14316_/A VGND VGND VPWR VPWR _14316_/X sky130_fd_sc_hd__buf_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18084_ _18008_/A VGND VGND VPWR VPWR _18084_/X sky130_fd_sc_hd__buf_2
X_15296_ _25013_/Q _15357_/A VGND VGND VPWR VPWR _15297_/C sky130_fd_sc_hd__or2_4
X_17035_ _24404_/Q VGND VGND VPWR VPWR _17035_/Y sky130_fd_sc_hd__inv_2
X_14247_ _25200_/Q VGND VGND VPWR VPWR _14247_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20416__A3 _20249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14178_ _25137_/Q VGND VGND VPWR VPWR _14178_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12592__A2_N _24864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _20789_/A _20790_/B _13129_/C _13128_/X VGND VGND VPWR VPWR _20794_/B sky130_fd_sc_hd__or4_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18986_ _14674_/A VGND VGND VPWR VPWR _18986_/X sky130_fd_sc_hd__buf_2
XANTENNA__24882__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14500__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21375__A _21375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17937_ _17929_/A _17924_/Y _17933_/X VGND VGND VPWR VPWR _17937_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24811__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17868_ _17868_/A VGND VGND VPWR VPWR _24273_/D sky130_fd_sc_hd__inv_2
XFILLER_27_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16253__B1 _16252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19605_/Y _19601_/X _19421_/X _19606_/X VGND VGND VPWR VPWR _23690_/D sky130_fd_sc_hd__a2bb2o_4
X_16819_ _16818_/Y _16816_/X _15734_/X _16816_/X VGND VGND VPWR VPWR _16819_/X sky130_fd_sc_hd__a2bb2o_4
X_17799_ _17771_/X _17780_/X _17750_/Y VGND VGND VPWR VPWR _17799_/X sky130_fd_sc_hd__o21a_4
XFILLER_242_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19538_ _19538_/A VGND VGND VPWR VPWR _21826_/B sky130_fd_sc_hd__inv_2
X_19469_ _19468_/Y _19466_/X _19377_/X _19466_/X VGND VGND VPWR VPWR _19469_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21500_ _21493_/X _21498_/X _21499_/X VGND VGND VPWR VPWR _21500_/X sky130_fd_sc_hd__o21a_4
XFILLER_195_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13621__A _18023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22480_ _22480_/A _22472_/Y _22480_/C _22480_/D VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__or4_4
XANTENNA__22934__A _22934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21431_ _21430_/X VGND VGND VPWR VPWR _21431_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_107_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24020_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_194_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24150_ _24145_/CLK _18762_/X HRESETn VGND VGND VPWR VPWR _24150_/Q sky130_fd_sc_hd__dfrtp_4
X_21362_ SSn_S3 _12108_/B SSn_S2 _13504_/B VGND VGND VPWR VPWR _21362_/X sky130_fd_sc_hd__o22a_4
X_20313_ _20312_/Y _20308_/X _20003_/X _20308_/X VGND VGND VPWR VPWR _23439_/D sky130_fd_sc_hd__a2bb2o_4
X_23101_ _15051_/A _22968_/B _22853_/X VGND VGND VPWR VPWR _23101_/X sky130_fd_sc_hd__and3_4
X_24081_ _25365_/CLK _20437_/A HRESETn VGND VGND VPWR VPWR _15493_/A sky130_fd_sc_hd__dfrtp_4
X_21293_ _21121_/X VGND VGND VPWR VPWR _21293_/X sky130_fd_sc_hd__buf_2
XFILLER_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23032_ _13659_/C _21306_/A _13129_/C _21607_/X VGND VGND VPWR VPWR _23032_/Y sky130_fd_sc_hd__a22oi_4
X_20244_ _20242_/Y _20240_/X _20243_/X _20240_/X VGND VGND VPWR VPWR _23465_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15819__B1 _11787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16087__A3 _15933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20175_ _20174_/Y _20172_/X _20105_/X _20172_/X VGND VGND VPWR VPWR _20175_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21285__A _25062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15834__A3 _16252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24983_ _24981_/CLK _15429_/X HRESETn VGND VGND VPWR VPWR _24983_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24552__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16379__A _16379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23934_ _24111_/CLK _23934_/D VGND VGND VPWR VPWR _23934_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23865_ _23577_/CLK _23865_/D VGND VGND VPWR VPWR _23865_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22816_ _23148_/A VGND VGND VPWR VPWR _22816_/X sky130_fd_sc_hd__buf_2
X_23796_ _24214_/CLK _23796_/D VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_232_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25535_ _25539_/CLK _25535_/D HRESETn VGND VGND VPWR VPWR _25535_/Q sky130_fd_sc_hd__dfrtp_4
X_22747_ _24062_/Q _21320_/A _13142_/C _21322_/X VGND VGND VPWR VPWR _22747_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_197_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12500_ _12278_/Y _12500_/B VGND VGND VPWR VPWR _12500_/Y sky130_fd_sc_hd__nand2_4
X_13480_ _13480_/A VGND VGND VPWR VPWR _13480_/Y sky130_fd_sc_hd__inv_2
X_25466_ _25456_/CLK _12413_/Y HRESETn VGND VGND VPWR VPWR _25466_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_66_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_66_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22678_ _22678_/A _22678_/B VGND VGND VPWR VPWR _22678_/X sky130_fd_sc_hd__or2_4
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22844__A _23087_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12431_ _12430_/X VGND VGND VPWR VPWR _12431_/Y sky130_fd_sc_hd__inv_2
X_24417_ _24684_/CLK _16873_/X HRESETn VGND VGND VPWR VPWR _20105_/A sky130_fd_sc_hd__dfrtp_4
X_21629_ _21629_/A _21629_/B VGND VGND VPWR VPWR _21629_/X sky130_fd_sc_hd__or2_4
XFILLER_138_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17938__A _13639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25397_ _24812_/CLK _12903_/Y HRESETn VGND VGND VPWR VPWR _25397_/Q sky130_fd_sc_hd__dfrtp_4
X_15150_ _15143_/X _15145_/X _15147_/X _15150_/D VGND VGND VPWR VPWR _15171_/B sky130_fd_sc_hd__or4_4
XFILLER_126_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12362_ _13006_/A _24838_/Q _13006_/A _24838_/Q VGND VGND VPWR VPWR _12362_/X sky130_fd_sc_hd__a2bb2o_4
X_24348_ _24354_/CLK _24348_/D HRESETn VGND VGND VPWR VPWR _24348_/Q sky130_fd_sc_hd__dfrtp_4
X_14101_ _14032_/A _20461_/C _14078_/X _14042_/B _14069_/B VGND VGND VPWR VPWR _25232_/D
+ sky130_fd_sc_hd__a32o_4
X_12293_ _12293_/A VGND VGND VPWR VPWR _12293_/Y sky130_fd_sc_hd__inv_2
X_15081_ _15196_/A _15193_/A VGND VGND VPWR VPWR _15081_/X sky130_fd_sc_hd__or2_4
X_24279_ _24283_/CLK _24279_/D HRESETn VGND VGND VPWR VPWR _17767_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14032_ _14032_/A _14032_/B VGND VGND VPWR VPWR _14054_/C sky130_fd_sc_hd__or2_4
XFILLER_180_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18840_ _18840_/A _18837_/X _18838_/X _18840_/D VGND VGND VPWR VPWR _18840_/X sky130_fd_sc_hd__or4_4
X_18771_ _18770_/X VGND VGND VPWR VPWR _24147_/D sky130_fd_sc_hd__inv_2
X_15983_ _15945_/Y VGND VGND VPWR VPWR _15983_/X sky130_fd_sc_hd__buf_2
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _21485_/A _17721_/X _21485_/A _17721_/X VGND VGND VPWR VPWR _17743_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14934_ _25032_/Q VGND VGND VPWR VPWR _15076_/C sky130_fd_sc_hd__inv_2
XANTENNA__12610__A _12609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17653_ _17578_/B _17649_/X VGND VGND VPWR VPWR _17653_/Y sky130_fd_sc_hd__nand2_4
X_14865_ _14837_/X _14864_/X _24962_/Q _14844_/X VGND VGND VPWR VPWR _14865_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16604_ _16618_/A VGND VGND VPWR VPWR _16604_/X sky130_fd_sc_hd__buf_2
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13816_ _13815_/Y _13813_/X _13524_/X _13813_/X VGND VGND VPWR VPWR _25277_/D sky130_fd_sc_hd__a2bb2o_4
X_17584_ _24307_/Q VGND VGND VPWR VPWR _17585_/C sky130_fd_sc_hd__inv_2
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14796_ _18059_/A VGND VGND VPWR VPWR _18027_/A sky130_fd_sc_hd__buf_2
XFILLER_235_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19323_ _19054_/A _19028_/B _19346_/C VGND VGND VPWR VPWR _19323_/X sky130_fd_sc_hd__or3_4
X_16535_ _16532_/Y _16533_/X _16534_/X _16533_/X VGND VGND VPWR VPWR _16535_/X sky130_fd_sc_hd__a2bb2o_4
X_13747_ _13747_/A VGND VGND VPWR VPWR _14772_/A sky130_fd_sc_hd__inv_2
XANTENNA__25428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19254_ _19139_/A VGND VGND VPWR VPWR _19254_/X sky130_fd_sc_hd__buf_2
XFILLER_231_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16466_ _16466_/A VGND VGND VPWR VPWR _16466_/Y sky130_fd_sc_hd__inv_2
X_13678_ _20831_/B VGND VGND VPWR VPWR _20834_/B sky130_fd_sc_hd__inv_2
X_18205_ _17973_/A _18204_/X _24248_/Q _18031_/A VGND VGND VPWR VPWR _24248_/D sky130_fd_sc_hd__o22a_4
X_15417_ _15401_/B _15417_/B _15427_/C VGND VGND VPWR VPWR _24987_/D sky130_fd_sc_hd__and3_4
X_12629_ _12660_/A _12588_/Y _12629_/C _12628_/X VGND VGND VPWR VPWR _12630_/B sky130_fd_sc_hd__or4_4
X_19185_ _19183_/Y _19181_/X _19184_/X _19181_/X VGND VGND VPWR VPWR _19185_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16397_ _24611_/Q VGND VGND VPWR VPWR _16397_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12057__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16752__A _16762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18136_ _18168_/A _18136_/B VGND VGND VPWR VPWR _18136_/X sky130_fd_sc_hd__or2_4
X_15348_ _15357_/A VGND VGND VPWR VPWR _15348_/X sky130_fd_sc_hd__buf_2
XANTENNA__25010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18067_ _13625_/X _18067_/B _18067_/C VGND VGND VPWR VPWR _18068_/C sky130_fd_sc_hd__and3_4
XFILLER_208_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15279_ _15276_/A _15276_/B VGND VGND VPWR VPWR _15279_/Y sky130_fd_sc_hd__nand2_4
XFILLER_160_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17018_ _17018_/A VGND VGND VPWR VPWR _17057_/B sky130_fd_sc_hd__inv_2
XFILLER_144_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22795__B1 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23339__A2 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15816__A3 _15738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18969_ _19085_/A VGND VGND VPWR VPWR _18969_/X sky130_fd_sc_hd__buf_2
XFILLER_227_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21980_ _14635_/Y _19610_/X VGND VGND VPWR VPWR _21980_/X sky130_fd_sc_hd__and2_4
XFILLER_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22929__A _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20931_ _20904_/A VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__buf_2
XPHY_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20862_ _20861_/X VGND VGND VPWR VPWR _24053_/D sky130_fd_sc_hd__inv_2
X_23650_ _23644_/CLK _19726_/X VGND VGND VPWR VPWR _13295_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22601_ _24663_/Q _16382_/A VGND VGND VPWR VPWR _22601_/X sky130_fd_sc_hd__or2_4
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20793_ _20788_/X _20791_/X _15594_/A _20792_/X VGND VGND VPWR VPWR _20793_/X sky130_fd_sc_hd__a2bb2o_4
X_23581_ _24217_/CLK _19922_/X VGND VGND VPWR VPWR _19921_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25320_ _25316_/CLK _13509_/X HRESETn VGND VGND VPWR VPWR _25320_/Q sky130_fd_sc_hd__dfrtp_4
X_22532_ _22296_/X _22530_/X _21124_/X _22531_/X VGND VGND VPWR VPWR _22535_/A sky130_fd_sc_hd__o22a_4
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25251_ _25253_/CLK _25251_/D HRESETn VGND VGND VPWR VPWR _21568_/A sky130_fd_sc_hd__dfrtp_4
X_22463_ _16527_/Y _21085_/X _16468_/A _16612_/Y _16552_/A VGND VGND VPWR VPWR _22463_/X
+ sky130_fd_sc_hd__o32a_4
X_24202_ _24201_/CLK _24202_/D HRESETn VGND VGND VPWR VPWR _24202_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21286__B1 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21414_ _21398_/X _21414_/B VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__or2_4
X_22394_ _22394_/A _20190_/Y VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__or2_4
X_25182_ _24112_/CLK _14321_/X HRESETn VGND VGND VPWR VPWR _25182_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11774__B1 _11773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21345_ _24553_/Q _22610_/B _21344_/X VGND VGND VPWR VPWR _21345_/X sky130_fd_sc_hd__o21a_4
X_24133_ _24138_/CLK _24133_/D HRESETn VGND VGND VPWR VPWR _24133_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21276_ _21272_/X _21275_/X _14692_/A VGND VGND VPWR VPWR _21277_/C sky130_fd_sc_hd__o21a_4
X_24064_ _24431_/CLK _20913_/X HRESETn VGND VGND VPWR VPWR _24064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12414__B _13017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24733__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_8_0_HCLK clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20227_ _21622_/B _20226_/X _16887_/X _20226_/X VGND VGND VPWR VPWR _23471_/D sky130_fd_sc_hd__a2bb2o_4
X_23015_ _21331_/X VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__buf_2
XANTENNA__22830__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16465__B1 _16375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20158_ _23497_/Q VGND VGND VPWR VPWR _21924_/B sky130_fd_sc_hd__inv_2
XFILLER_218_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19403__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12980_ _12796_/Y _12986_/B VGND VGND VPWR VPWR _12984_/B sky130_fd_sc_hd__or2_4
X_20089_ _20088_/Y _20086_/X _19728_/X _20086_/X VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__a2bb2o_4
X_24966_ _24966_/CLK _15467_/X HRESETn VGND VGND VPWR VPWR _13936_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__14727__A1_N _14725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22839__A _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11931_ _19990_/A VGND VGND VPWR VPWR _19626_/A sky130_fd_sc_hd__buf_2
X_23917_ _23918_/CLK _18957_/X VGND VGND VPWR VPWR _23917_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24897_ _24913_/CLK _24897_/D HRESETn VGND VGND VPWR VPWR _21026_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_57_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14650_ _17941_/A _17950_/A _14650_/C _18016_/A VGND VGND VPWR VPWR _14650_/X sky130_fd_sc_hd__and4_4
X_11862_ _14412_/A VGND VGND VPWR VPWR _11862_/X sky130_fd_sc_hd__buf_2
X_23848_ _24100_/CLK _23848_/D VGND VGND VPWR VPWR _23848_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13601_/A _13601_/B VGND VGND VPWR VPWR _13643_/A sky130_fd_sc_hd__or2_4
XFILLER_233_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14581_/A _14580_/Y VGND VGND VPWR VPWR _14582_/A sky130_fd_sc_hd__or2_4
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ HWDATA[19] VGND VGND VPWR VPWR _11793_/X sky130_fd_sc_hd__buf_2
X_23779_ _23850_/CLK _19351_/X VGND VGND VPWR VPWR _18012_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22710__B1 _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _16325_/A VGND VGND VPWR VPWR _16320_/X sky130_fd_sc_hd__buf_2
XANTENNA__13261__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _25188_/Q _13532_/B VGND VGND VPWR VPWR _13532_/X sky130_fd_sc_hd__or2_4
X_25518_ _23678_/CLK _25518_/D HRESETn VGND VGND VPWR VPWR _11886_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22574__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16251_ _16264_/A VGND VGND VPWR VPWR _16251_/X sky130_fd_sc_hd__buf_2
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13463_ _13315_/A _13459_/X _13462_/X VGND VGND VPWR VPWR _13463_/X sky130_fd_sc_hd__or3_4
X_25449_ _25454_/CLK _25449_/D HRESETn VGND VGND VPWR VPWR _25449_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15202_ _15079_/A _15201_/X VGND VGND VPWR VPWR _15202_/X sky130_fd_sc_hd__or2_4
X_12414_ _12414_/A _13017_/B VGND VGND VPWR VPWR _12414_/X sky130_fd_sc_hd__or2_4
XFILLER_145_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16182_ _14778_/X _16182_/B VGND VGND VPWR VPWR _16182_/X sky130_fd_sc_hd__and2_4
X_13394_ _13282_/A _19710_/A VGND VGND VPWR VPWR _13394_/X sky130_fd_sc_hd__or2_4
XFILLER_138_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_153_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25188_/CLK sky130_fd_sc_hd__clkbuf_1
X_15133_ _24998_/Q _15131_/Y _15399_/A _15135_/A VGND VGND VPWR VPWR _15133_/X sky130_fd_sc_hd__a2bb2o_4
X_12345_ _25358_/Q VGND VGND VPWR VPWR _13068_/A sky130_fd_sc_hd__inv_2
XFILLER_181_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15064_ _15064_/A _15064_/B _15056_/X _15063_/X VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__or4_4
X_19941_ _19940_/Y _19938_/X _19810_/X _19938_/X VGND VGND VPWR VPWR _19941_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12276_ _12275_/Y _24783_/Q _12275_/Y _24783_/Q VGND VGND VPWR VPWR _12280_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14015_ _14058_/A _14015_/B _13999_/D _14015_/D VGND VGND VPWR VPWR _14552_/A sky130_fd_sc_hd__and4_4
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19872_ _21782_/B _19867_/X _19803_/X _19867_/X VGND VGND VPWR VPWR _23600_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18823_ _18689_/A _18825_/B _18822_/Y VGND VGND VPWR VPWR _24134_/D sky130_fd_sc_hd__o21a_4
XFILLER_110_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15966_ _12266_/Y _15962_/X _15965_/X _15962_/X VGND VGND VPWR VPWR _24773_/D sky130_fd_sc_hd__a2bb2o_4
X_18754_ _18756_/B VGND VGND VPWR VPWR _18755_/B sky130_fd_sc_hd__inv_2
XANTENNA__12340__A _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16208__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14917_ _14916_/Y VGND VGND VPWR VPWR _15256_/A sky130_fd_sc_hd__buf_2
X_17705_ _17671_/X VGND VGND VPWR VPWR _17705_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15897_ _15894_/X _15895_/X _15748_/X _24806_/Q _15896_/X VGND VGND VPWR VPWR _15897_/X
+ sky130_fd_sc_hd__a32o_4
X_18685_ _24135_/Q VGND VGND VPWR VPWR _18685_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15651__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14848_ _14848_/A VGND VGND VPWR VPWR _14848_/Y sky130_fd_sc_hd__inv_2
X_17636_ _17579_/C _17635_/X VGND VGND VPWR VPWR _17636_/X sky130_fd_sc_hd__or2_4
XFILLER_208_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12577__A1_N _12618_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17567_ _24719_/Q VGND VGND VPWR VPWR _17567_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14779_ _14779_/A _14769_/X _13599_/B VGND VGND VPWR VPWR _14790_/B sky130_fd_sc_hd__and3_4
XFILLER_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17708__B1 _17611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__B2 _22644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13171__A _13423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16518_ _16517_/Y _16513_/X _16248_/X _16513_/X VGND VGND VPWR VPWR _24564_/D sky130_fd_sc_hd__a2bb2o_4
X_19306_ _19304_/Y _19302_/X _19305_/X _19302_/X VGND VGND VPWR VPWR _19306_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17498_ _13183_/X _17497_/Y _13171_/X _17496_/X VGND VGND VPWR VPWR _17498_/X sky130_fd_sc_hd__o22a_4
XFILLER_210_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22484__A _22157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16449_ _16448_/Y _16446_/X _16368_/X _16446_/X VGND VGND VPWR VPWR _16449_/X sky130_fd_sc_hd__a2bb2o_4
X_19237_ _19232_/Y _19236_/X _19169_/X _19236_/X VGND VGND VPWR VPWR _23820_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16482__A _16482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19168_ _19181_/A VGND VGND VPWR VPWR _19168_/X sky130_fd_sc_hd__buf_2
XFILLER_145_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11756__B1 _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18119_ _14656_/A _18119_/B _18118_/X VGND VGND VPWR VPWR _18119_/X sky130_fd_sc_hd__and3_4
XFILLER_191_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19099_ _19099_/A VGND VGND VPWR VPWR _19099_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12515__A _13017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21130_ _21130_/A _21046_/X VGND VGND VPWR VPWR _21130_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16695__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21828__A _21668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21061_ _11728_/X VGND VGND VPWR VPWR _21062_/A sky130_fd_sc_hd__inv_2
XANTENNA__15826__A _15826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20012_ _20012_/A VGND VGND VPWR VPWR _21187_/B sky130_fd_sc_hd__inv_2
XANTENNA__16447__B1 _16364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24820_ _24856_/CLK _24820_/D HRESETn VGND VGND VPWR VPWR _23290_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24751_ _24735_/CLK _24751_/D HRESETn VGND VGND VPWR VPWR _16008_/A sky130_fd_sc_hd__dfrtp_4
X_21963_ _21948_/A _19635_/Y VGND VGND VPWR VPWR _21964_/C sky130_fd_sc_hd__or2_4
X_23702_ _23669_/CLK _23702_/D VGND VGND VPWR VPWR _19568_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_214_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20914_ _20915_/B VGND VGND VPWR VPWR _20914_/Y sky130_fd_sc_hd__inv_2
XFILLER_242_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24682_ _24169_/CLK _24682_/D HRESETn VGND VGND VPWR VPWR _23309_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21894_ _21914_/A _21894_/B VGND VGND VPWR VPWR _21894_/X sky130_fd_sc_hd__or2_4
XFILLER_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23644_/CLK _19776_/X VGND VGND VPWR VPWR _23633_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A VGND VGND VPWR VPWR _20845_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _23513_/CLK _23564_/D VGND VGND VPWR VPWR _19964_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ _20776_/A _24033_/Q _20768_/A _20768_/B VGND VGND VPWR VPWR _20776_/X sky130_fd_sc_hd__or4_4
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25303_ _25188_/CLK _13683_/X HRESETn VGND VGND VPWR VPWR _25303_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22515_ _22459_/X _22512_/X _22462_/X _22514_/X VGND VGND VPWR VPWR _22516_/B sky130_fd_sc_hd__o22a_4
XFILLER_167_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _23494_/CLK _23495_/D VGND VGND VPWR VPWR _23495_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25234_ _25105_/CLK _14097_/X HRESETn VGND VGND VPWR VPWR _13994_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22446_ _22446_/A _22445_/X VGND VGND VPWR VPWR _22446_/Y sky130_fd_sc_hd__nor2_4
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24914__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25165_ _24121_/CLK _14370_/X HRESETn VGND VGND VPWR VPWR _25165_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22377_ _22373_/X _22376_/X _21785_/X VGND VGND VPWR VPWR _22377_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_226_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _25125_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14651__A1_N _18069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12130_ _25475_/Q VGND VGND VPWR VPWR _12175_/A sky130_fd_sc_hd__inv_2
X_24116_ _24119_/CLK _20981_/X HRESETn VGND VGND VPWR VPWR _12136_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16686__B1 _16417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21328_ _21874_/A VGND VGND VPWR VPWR _22945_/A sky130_fd_sc_hd__buf_2
X_25096_ _25093_/CLK _14604_/X HRESETn VGND VGND VPWR VPWR _25096_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22759__B1 _24840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12061_ _12061_/A _12061_/B VGND VGND VPWR VPWR _13476_/D sky130_fd_sc_hd__or2_4
X_21259_ _21259_/A _20145_/Y VGND VGND VPWR VPWR _21260_/C sky130_fd_sc_hd__or2_4
X_24047_ _24485_/CLK _20838_/Y HRESETn VGND VGND VPWR VPWR _24047_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15820_ _12375_/Y _15818_/X _11790_/X _15818_/X VGND VGND VPWR VPWR _24845_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12376__A2_N _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22569__A _21129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15751_ _15751_/A VGND VGND VPWR VPWR _15751_/X sky130_fd_sc_hd__buf_2
XANTENNA__21473__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12963_ _12793_/A _12962_/Y VGND VGND VPWR VPWR _12963_/X sky130_fd_sc_hd__or2_4
X_24949_ _23717_/CLK _15509_/X HRESETn VGND VGND VPWR VPWR _11736_/A sky130_fd_sc_hd__dfrtp_4
X_14702_ _22228_/A VGND VGND VPWR VPWR _21630_/A sky130_fd_sc_hd__buf_2
X_11914_ _11905_/X _11908_/Y _11913_/Y VGND VGND VPWR VPWR _11914_/X sky130_fd_sc_hd__o21a_4
X_18470_ _24177_/Q VGND VGND VPWR VPWR _18471_/D sky130_fd_sc_hd__inv_2
X_15682_ _15681_/X VGND VGND VPWR VPWR _16382_/A sky130_fd_sc_hd__buf_2
X_12894_ _12894_/A VGND VGND VPWR VPWR _25399_/D sky130_fd_sc_hd__inv_2
XFILLER_245_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17421_ _14816_/A VGND VGND VPWR VPWR _20680_/A sky130_fd_sc_hd__buf_2
X_14633_ _25086_/Q _13645_/X _14632_/X VGND VGND VPWR VPWR _14633_/X sky130_fd_sc_hd__a21o_4
X_11845_ _11803_/X VGND VGND VPWR VPWR _11845_/X sky130_fd_sc_hd__buf_2
XFILLER_233_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17351_/X VGND VGND VPWR VPWR _17352_/Y sky130_fd_sc_hd__inv_2
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14611_/A _13599_/B VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__or2_4
XFILLER_186_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ HWDATA[24] VGND VGND VPWR VPWR _11776_/X sky130_fd_sc_hd__buf_2
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16302_/Y _16298_/X _15952_/X _16298_/X VGND VGND VPWR VPWR _24644_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13515_ _13514_/Y _13510_/X _11851_/X _13510_/X VGND VGND VPWR VPWR _25317_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17283_ _17243_/X _17283_/B VGND VGND VPWR VPWR _17286_/B sky130_fd_sc_hd__or2_4
XFILLER_13_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14495_ _21726_/A _14490_/X _14412_/X _14490_/X VGND VGND VPWR VPWR _14495_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_36_0_HCLK clkbuf_6_36_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _19022_/A VGND VGND VPWR VPWR _19022_/Y sky130_fd_sc_hd__inv_2
X_16234_ _16202_/A VGND VGND VPWR VPWR _16264_/A sky130_fd_sc_hd__buf_2
X_13446_ _13317_/A _13446_/B VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__or2_4
XFILLER_167_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24655__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16165_ _16164_/Y _16162_/X _16073_/X _16162_/X VGND VGND VPWR VPWR _16165_/X sky130_fd_sc_hd__a2bb2o_4
X_13377_ _13207_/X _13376_/X _25334_/Q _13267_/X VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__o22a_4
XFILLER_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22751__B _22589_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15116_ _15116_/A _15116_/B _15112_/X _15116_/D VGND VGND VPWR VPWR _15116_/X sky130_fd_sc_hd__or4_4
XFILLER_154_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12328_ _25348_/Q _12327_/A _12326_/Y _12327_/Y VGND VGND VPWR VPWR _12335_/B sky130_fd_sc_hd__o22a_4
XFILLER_142_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16096_ _16096_/A VGND VGND VPWR VPWR _16096_/X sky130_fd_sc_hd__buf_2
XFILLER_108_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15047_ _14956_/Y VGND VGND VPWR VPWR _15248_/A sky130_fd_sc_hd__buf_2
X_19924_ _18914_/A _13761_/X _13762_/X _13770_/X VGND VGND VPWR VPWR _19925_/A sky130_fd_sc_hd__or4_4
X_12259_ _12464_/A _22758_/A _12464_/A _22758_/A VGND VGND VPWR VPWR _12259_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14550__A _14550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16429__B1 _16241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19855_ _23605_/Q VGND VGND VPWR VPWR _21241_/B sky130_fd_sc_hd__inv_2
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18806_ _18806_/A _18806_/B _18805_/X VGND VGND VPWR VPWR _18806_/X sky130_fd_sc_hd__and3_4
XFILLER_228_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13166__A _13451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19786_ _23628_/Q VGND VGND VPWR VPWR _19786_/Y sky130_fd_sc_hd__inv_2
X_16998_ _16998_/A _16993_/X _16995_/X _16998_/D VGND VGND VPWR VPWR _16998_/X sky130_fd_sc_hd__or4_4
XFILLER_205_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22479__A _22479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23175__B1 _25399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18737_ _18737_/A _18736_/Y VGND VGND VPWR VPWR _18739_/B sky130_fd_sc_hd__or2_4
XFILLER_95_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12466__A1 _12247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15949_ _12226_/Y _15947_/X _15948_/X _15947_/X VGND VGND VPWR VPWR _24782_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_243_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21725__A1 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18668_ _16625_/Y _24134_/Q _24521_/Q _18689_/C VGND VGND VPWR VPWR _18673_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17619_ _17895_/B _17615_/B _17618_/X VGND VGND VPWR VPWR _17620_/A sky130_fd_sc_hd__or3_4
XFILLER_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_237_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18599_ _18565_/X VGND VGND VPWR VPWR _18599_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20630_ _15482_/Y _20623_/X _20680_/A _20629_/X VGND VGND VPWR VPWR _20631_/A sky130_fd_sc_hd__a211o_4
XFILLER_32_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20561_ _18878_/X _20561_/B _20556_/X VGND VGND VPWR VPWR _20561_/X sky130_fd_sc_hd__and3_4
XANTENNA__23103__A _21879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22300_ _22296_/X _22297_/X _22298_/X _22299_/X VGND VGND VPWR VPWR _22301_/B sky130_fd_sc_hd__o22a_4
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20492_ _15465_/A _20682_/B _20487_/B VGND VGND VPWR VPWR _20537_/A sky130_fd_sc_hd__and3_4
X_23280_ _23280_/A _23279_/X VGND VGND VPWR VPWR _23280_/Y sky130_fd_sc_hd__nor2_4
XFILLER_118_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22231_ _22227_/A _19261_/Y VGND VGND VPWR VPWR _22231_/X sky130_fd_sc_hd__or2_4
XFILLER_192_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16668__B1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22162_ _22162_/A _22155_/B VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__or2_4
XFILLER_172_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21113_ _21064_/X VGND VGND VPWR VPWR _21113_/X sky130_fd_sc_hd__buf_2
XFILLER_246_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15556__A _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22093_ _22093_/A _20176_/Y VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_56_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _24238_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21044_ _24790_/Q _21069_/B VGND VGND VPWR VPWR _21044_/X sky130_fd_sc_hd__or2_4
XANTENNA__22756__A3 _22303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22389__A _22090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24956__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24803_ _24803_/CLK _15900_/X HRESETn VGND VGND VPWR VPWR _22669_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16840__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22995_ _22993_/X _22994_/X _22503_/X _25546_/Q _22793_/X VGND VGND VPWR VPWR _22995_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_228_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21716__A1 _15565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21724__C _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21716__B2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24734_ _24735_/CLK _24734_/D HRESETn VGND VGND VPWR VPWR _16051_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13804__A _16464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21946_ _21936_/A VGND VGND VPWR VPWR _21947_/A sky130_fd_sc_hd__buf_2
XANTENNA__25113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24665_ _24674_/CLK _16246_/X HRESETn VGND VGND VPWR VPWR _16244_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _15036_/A _21877_/B _21096_/X VGND VGND VPWR VPWR _21877_/X sky130_fd_sc_hd__and3_4
XFILLER_242_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _25507_/CLK _23616_/D VGND VGND VPWR VPWR _23616_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20698_/X _20827_/X _24928_/Q _20744_/A VGND VGND VPWR VPWR _20828_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24596_ _24592_/CLK _24596_/D HRESETn VGND VGND VPWR VPWR _16434_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_202_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18345__B1 _17485_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23547_ _23563_/CLK _23547_/D VGND VGND VPWR VPWR _23547_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20759_ _20756_/Y _20757_/Y _20758_/X VGND VGND VPWR VPWR _20759_/X sky130_fd_sc_hd__o21a_4
XFILLER_11_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22692__A2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13372_/A _19821_/A VGND VGND VPWR VPWR _13301_/C sky130_fd_sc_hd__or2_4
XFILLER_11_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _14268_/A VGND VGND VPWR VPWR _14280_/X sky130_fd_sc_hd__buf_2
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23478_ _23494_/CLK _23478_/D VGND VGND VPWR VPWR _23478_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ _13317_/A _18963_/A VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__or2_4
X_25217_ _25215_/CLK _14185_/Y HRESETn VGND VGND VPWR VPWR _14174_/A sky130_fd_sc_hd__dfrtp_4
X_22429_ _21431_/X _22428_/X _22303_/X _24867_/Q _22558_/A VGND VGND VPWR VPWR _22430_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22571__B _22610_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13162_ _13192_/A _13162_/B VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__or2_4
X_25148_ _25148_/CLK _14429_/X HRESETn VGND VGND VPWR VPWR _14425_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__21652__B1 _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21468__A _22271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12113_ _25482_/Q VGND VGND VPWR VPWR _12113_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13093_ _12332_/Y _13092_/X VGND VGND VPWR VPWR _13106_/B sky130_fd_sc_hd__or2_4
X_17970_ _15686_/X _15693_/A _14628_/Y _15926_/X VGND VGND VPWR VPWR _17973_/A sky130_fd_sc_hd__a211o_4
X_25079_ _23836_/CLK _25079_/D HRESETn VGND VGND VPWR VPWR _25079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12044_ _12042_/Y _12038_/X _25497_/Q _12043_/X VGND VGND VPWR VPWR _25498_/D sky130_fd_sc_hd__a2bb2o_4
X_16921_ _22413_/A _24270_/Q _16159_/Y _16920_/Y VGND VGND VPWR VPWR _16921_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19640_ _19638_/Y _19633_/X _19639_/X _19633_/X VGND VGND VPWR VPWR _19640_/X sky130_fd_sc_hd__a2bb2o_4
X_16852_ _14931_/Y _16849_/X _16530_/X _16849_/X VGND VGND VPWR VPWR _24426_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16831__B1 HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15803_ _15790_/X _15797_/X _15562_/X _24856_/Q _15802_/X VGND VGND VPWR VPWR _24856_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_207_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16783_ _15022_/Y _16779_/X _16609_/X _16782_/X VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__a2bb2o_4
X_19571_ _19570_/Y _19565_/X _19410_/X _19565_/A VGND VGND VPWR VPWR _23701_/D sky130_fd_sc_hd__a2bb2o_4
X_13995_ _14032_/B VGND VGND VPWR VPWR _14004_/A sky130_fd_sc_hd__inv_2
XFILLER_206_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16297__A _16290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22904__B1 _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15734_ HWDATA[25] VGND VGND VPWR VPWR _15734_/X sky130_fd_sc_hd__buf_2
X_18522_ _18516_/B VGND VGND VPWR VPWR _18523_/B sky130_fd_sc_hd__inv_2
X_12946_ _12941_/A _12940_/X _12891_/X _12942_/Y VGND VGND VPWR VPWR _12947_/A sky130_fd_sc_hd__a211o_4
XFILLER_246_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17387__A1 _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15665_ _15661_/X VGND VGND VPWR VPWR _21105_/B sky130_fd_sc_hd__buf_2
X_18453_ _16199_/Y _24193_/Q _16199_/Y _24193_/Q VGND VGND VPWR VPWR _18453_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12877_ _12876_/X VGND VGND VPWR VPWR _25403_/D sky130_fd_sc_hd__inv_2
XFILLER_221_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15937__A2 _15796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14613_/B _14615_/Y _14608_/X _14611_/X _13582_/A VGND VGND VPWR VPWR _14616_/X
+ sky130_fd_sc_hd__a32o_4
X_17404_ _17404_/A _17404_/B VGND VGND VPWR VPWR _20661_/A sky130_fd_sc_hd__or2_4
XPHY_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11824_/Y _11825_/X _11827_/X _11825_/X VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__a2bb2o_4
X_18384_ _18379_/A VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__buf_2
XFILLER_178_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15596_ _24918_/Q VGND VGND VPWR VPWR _15596_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24836__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17335_ _17315_/X _17330_/X _17334_/X VGND VGND VPWR VPWR _24363_/D sky130_fd_sc_hd__and3_4
XFILLER_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14554_/A _14059_/B _14546_/X _14023_/X VGND VGND VPWR VPWR _14548_/A sky130_fd_sc_hd__or4_4
X_11759_ _11749_/X VGND VGND VPWR VPWR _11759_/X sky130_fd_sc_hd__buf_2
XANTENNA__22683__A2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18017__A _18097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17266_ _17266_/A _17231_/Y _17248_/X _17265_/X VGND VGND VPWR VPWR _17267_/B sky130_fd_sc_hd__or4_4
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14478_ HWDATA[1] VGND VGND VPWR VPWR _14479_/A sky130_fd_sc_hd__buf_2
XFILLER_186_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16217_ _23076_/A VGND VGND VPWR VPWR _16217_/Y sky130_fd_sc_hd__inv_2
X_19005_ _19001_/Y _19004_/X _17427_/X _19004_/X VGND VGND VPWR VPWR _23900_/D sky130_fd_sc_hd__a2bb2o_4
X_13429_ _13257_/X _13429_/B VGND VGND VPWR VPWR _13429_/X sky130_fd_sc_hd__or2_4
X_17197_ _24353_/Q VGND VGND VPWR VPWR _17197_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16148_ _16162_/A VGND VGND VPWR VPWR _16148_/X sky130_fd_sc_hd__buf_2
XANTENNA__21643__B1 _14721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21378__A _21565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16079_ _16078_/Y _16076_/X _15483_/X _16076_/X VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21528__D _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19907_ _19907_/A VGND VGND VPWR VPWR _22255_/B sky130_fd_sc_hd__inv_2
X_19838_ _19838_/A VGND VGND VPWR VPWR _19838_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19769_ HWDATA[6] VGND VGND VPWR VPWR _19769_/X sky130_fd_sc_hd__buf_2
XFILLER_244_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22002__A _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12206__A2_N _21091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21800_ _21660_/X _21798_/X _21519_/X _21799_/X VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__a211o_4
X_22780_ _22777_/X _22778_/X _22484_/X _24841_/Q _22779_/X VGND VGND VPWR VPWR _22780_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21731_ _21731_/A _21731_/B VGND VGND VPWR VPWR _21731_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20921__A2 _20854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24450_ _24473_/CLK _24450_/D HRESETn VGND VGND VPWR VPWR _16803_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21662_ _18278_/X _21659_/X _21519_/X _21661_/Y VGND VGND VPWR VPWR _21662_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23320__B1 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24577__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23401_ _23493_/CLK _23401_/D VGND VGND VPWR VPWR _23401_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20613_ _20613_/A VGND VGND VPWR VPWR _20613_/Y sky130_fd_sc_hd__inv_2
X_24381_ _24383_/CLK _17167_/X HRESETn VGND VGND VPWR VPWR _24381_/Q sky130_fd_sc_hd__dfrtp_4
X_21593_ _16544_/Y _21752_/B VGND VGND VPWR VPWR _21593_/X sky130_fd_sc_hd__and2_4
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16064__A1_N _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23332_ _23332_/A _21711_/A VGND VGND VPWR VPWR _23332_/X sky130_fd_sc_hd__and2_4
X_20544_ _20683_/A _20486_/Y _20501_/B _20543_/X VGND VGND VPWR VPWR _20544_/X sky130_fd_sc_hd__a211o_4
XFILLER_192_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22672__A _22155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23263_ _23025_/A _23260_/X _23263_/C VGND VGND VPWR VPWR _23263_/X sky130_fd_sc_hd__and3_4
XANTENNA__19827__B1 _19753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20475_ _20463_/A _20471_/B _20475_/C _20477_/C VGND VGND VPWR VPWR _20476_/D sky130_fd_sc_hd__and4_4
XFILLER_180_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25002_ _25002_/CLK _25002_/D HRESETn VGND VGND VPWR VPWR _25002_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22214_ _22214_/A _22214_/B _22214_/C VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__or3_4
XFILLER_146_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23194_ _23156_/A _23182_/Y _23187_/X _23194_/D VGND VGND VPWR VPWR _23194_/X sky130_fd_sc_hd__or4_4
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15286__A _15292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22145_ _21306_/A _22145_/B _22145_/C VGND VGND VPWR VPWR _22145_/X sky130_fd_sc_hd__and3_4
XFILLER_133_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22076_ _22071_/X _22075_/X _21785_/X VGND VGND VPWR VPWR _22076_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21027_ _15709_/X VGND VGND VPWR VPWR _21027_/X sky130_fd_sc_hd__buf_2
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16813__B1 HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23008__A _23008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12800_ _12800_/A _12772_/X _12800_/C _12799_/X VGND VGND VPWR VPWR _12846_/A sky130_fd_sc_hd__or4_4
X_13780_ _14684_/A VGND VGND VPWR VPWR _13781_/A sky130_fd_sc_hd__buf_2
XFILLER_90_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22978_ _22973_/Y _22977_/Y _22868_/X VGND VGND VPWR VPWR _22978_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12731_ _12731_/A _12729_/Y _12741_/C VGND VGND VPWR VPWR _25412_/D sky130_fd_sc_hd__and3_4
X_24717_ _24689_/CLK _16099_/X HRESETn VGND VGND VPWR VPWR _24717_/Q sky130_fd_sc_hd__dfrtp_4
X_21929_ _21913_/X _21928_/X _21288_/X VGND VGND VPWR VPWR _21929_/X sky130_fd_sc_hd__a21o_4
XFILLER_204_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20373__B1 _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15450_ _14255_/X _15447_/A VGND VGND VPWR VPWR _15450_/Y sky130_fd_sc_hd__nor2_4
X_12662_ _12640_/B VGND VGND VPWR VPWR _12662_/X sky130_fd_sc_hd__buf_2
X_24648_ _24641_/CLK _24648_/D HRESETn VGND VGND VPWR VPWR _24648_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_203_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _20514_/D _14391_/X _14400_/X _14393_/X VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23311__B1 _22852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15384_/A _15381_/B _15380_/Y VGND VGND VPWR VPWR _24997_/D sky130_fd_sc_hd__and3_4
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12593_/A VGND VGND VPWR VPWR _12593_/Y sky130_fd_sc_hd__inv_2
X_24579_ _24562_/CLK _24579_/D HRESETn VGND VGND VPWR VPWR _24579_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17042_/B _17120_/B VGND VGND VPWR VPWR _17120_/Y sky130_fd_sc_hd__nand2_4
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _25176_/Q _14320_/A _14316_/X _13502_/A _14315_/A VGND VGND VPWR VPWR _25176_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_21_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17051_ _17051_/A VGND VGND VPWR VPWR _17051_/Y sky130_fd_sc_hd__inv_2
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _25197_/Q VGND VGND VPWR VPWR _14263_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15552__B1 HADDR[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19818__B1 _19817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22417__A2 _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19594__C _13786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16002_ _16001_/X VGND VGND VPWR VPWR _16288_/B sky130_fd_sc_hd__inv_2
X_13214_ _13271_/A VGND VGND VPWR VPWR _13450_/A sky130_fd_sc_hd__buf_2
XFILLER_167_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14194_ _20511_/A VGND VGND VPWR VPWR _14194_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19294__B2 _19293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20187__A2_N _20184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13145_ _13145_/A _13145_/B _13145_/C _13144_/X VGND VGND VPWR VPWR _13145_/X sky130_fd_sc_hd__or4_4
XFILLER_151_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12613__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21926__A _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ _13069_/A _13066_/B _13075_/X VGND VGND VPWR VPWR _25355_/D sky130_fd_sc_hd__and3_4
X_17953_ _17949_/X _17952_/X _18016_/A VGND VGND VPWR VPWR _17954_/C sky130_fd_sc_hd__o21a_4
XFILLER_183_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12027_ _12023_/Y _20976_/A _12023_/Y _20976_/A VGND VGND VPWR VPWR _12027_/X sky130_fd_sc_hd__a2bb2o_4
X_16904_ _16899_/X _16904_/B _16904_/C _16904_/D VGND VGND VPWR VPWR _16932_/A sky130_fd_sc_hd__or4_4
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17884_ _17881_/A _17877_/B _17883_/X VGND VGND VPWR VPWR _24268_/D sky130_fd_sc_hd__and3_4
XANTENNA__18300__A _21212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19623_ _18282_/X _19480_/X _18289_/X VGND VGND VPWR VPWR _19623_/X sky130_fd_sc_hd__or3_4
X_16835_ _16832_/Y _16834_/X _15748_/X _16834_/X VGND VGND VPWR VPWR _24435_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13444__A _13153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19554_ _19554_/A VGND VGND VPWR VPWR _19554_/Y sky130_fd_sc_hd__inv_2
X_13978_ _13977_/Y _13978_/B VGND VGND VPWR VPWR _13978_/X sky130_fd_sc_hd__and2_4
X_16766_ _15039_/Y _16762_/X _16419_/X _16762_/X VGND VGND VPWR VPWR _24468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20125__A2_N _20118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18505_ _18828_/B VGND VGND VPWR VPWR _18505_/X sky130_fd_sc_hd__buf_2
XANTENNA__21661__A _13748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12929_ _12819_/A _12929_/B VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__or2_4
X_15717_ _22146_/B VGND VGND VPWR VPWR _15718_/A sky130_fd_sc_hd__buf_2
XFILLER_206_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16697_ _16685_/A VGND VGND VPWR VPWR _16697_/X sky130_fd_sc_hd__buf_2
X_19485_ _22357_/B _19484_/X _11939_/X _19484_/X VGND VGND VPWR VPWR _19485_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12841__B2 _24794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18436_ _16247_/Y _18475_/A _16247_/Y _18475_/A VGND VGND VPWR VPWR _18436_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19131__A _19131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15648_ _15647_/Y _15584_/A _15489_/X _15584_/A VGND VGND VPWR VPWR _24898_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24670__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15579_ _24925_/Q VGND VGND VPWR VPWR _23213_/A sky130_fd_sc_hd__inv_2
X_18367_ _18366_/Y _18361_/A _18366_/A _17492_/X VGND VGND VPWR VPWR _18368_/A sky130_fd_sc_hd__o22a_4
XFILLER_159_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17318_ _17318_/A _17326_/D VGND VGND VPWR VPWR _17318_/X sky130_fd_sc_hd__or2_4
XFILLER_187_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18298_ _24219_/Q VGND VGND VPWR VPWR _18301_/A sky130_fd_sc_hd__buf_2
XANTENNA__17532__A1 _25543_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17249_ _24357_/Q VGND VGND VPWR VPWR _17362_/A sky130_fd_sc_hd__inv_2
XFILLER_190_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15543__B1 HADDR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20260_ _20260_/A VGND VGND VPWR VPWR _20260_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20191_ _13774_/X _13761_/X _13762_/X _13770_/X VGND VGND VPWR VPWR _20191_/X sky130_fd_sc_hd__or4_4
XFILLER_227_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15846__A1 _15833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15809__A1_N _12337_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15846__B2 _15802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23950_ _23960_/CLK _20559_/Y HRESETn VGND VGND VPWR VPWR _20555_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22901_ _22171_/A VGND VGND VPWR VPWR _22950_/A sky130_fd_sc_hd__buf_2
XFILLER_243_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23881_ _23880_/CLK _23881_/D VGND VGND VPWR VPWR _23881_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22832_ _23025_/A _22832_/B _22831_/X VGND VGND VPWR VPWR _22832_/X sky130_fd_sc_hd__and3_4
XANTENNA__24758__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25551_ _24697_/CLK _11771_/X HRESETn VGND VGND VPWR VPWR _11768_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22763_ _22763_/A _23053_/A VGND VGND VPWR VPWR _22763_/X sky130_fd_sc_hd__or2_4
X_24502_ _24500_/CLK _24502_/D HRESETn VGND VGND VPWR VPWR _24502_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21714_ _21714_/A _21714_/B VGND VGND VPWR VPWR _21714_/X sky130_fd_sc_hd__and2_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21290__B _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25482_ _25316_/CLK _25482_/D HRESETn VGND VGND VPWR VPWR _25482_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22694_ _15613_/Y _22694_/B VGND VGND VPWR VPWR _22694_/X sky130_fd_sc_hd__and2_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24433_ _24431_/CLK _16840_/X HRESETn VGND VGND VPWR VPWR _24433_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21645_ _21783_/A _20071_/Y VGND VGND VPWR VPWR _21646_/C sky130_fd_sc_hd__or2_4
XANTENNA__22647__A2 _22646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24364_ _24629_/CLK _17332_/X HRESETn VGND VGND VPWR VPWR _24364_/Q sky130_fd_sc_hd__dfrtp_4
X_21576_ _21741_/A _21575_/X VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__and2_4
XANTENNA__17523__A1 _25532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23315_ _24449_/Q _22153_/X _22815_/X _23314_/X VGND VGND VPWR VPWR _23315_/X sky130_fd_sc_hd__a211o_4
X_20527_ _20527_/A _20526_/X VGND VGND VPWR VPWR _24089_/D sky130_fd_sc_hd__or2_4
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15534__B1 HADDR[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ _24295_/CLK _17746_/X HRESETn VGND VGND VPWR VPWR _21704_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23246_ _23137_/X _23244_/X _23139_/X _23245_/X VGND VGND VPWR VPWR _23247_/B sky130_fd_sc_hd__o22a_4
X_20458_ _20457_/X VGND VGND VPWR VPWR _20609_/B sky130_fd_sc_hd__buf_2
XFILLER_180_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19276__B2 _19258_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25307__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22280__B1 _21968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23177_ _16664_/Y _23177_/B VGND VGND VPWR VPWR _23177_/X sky130_fd_sc_hd__and2_4
X_20389_ _22252_/B _20386_/X _19629_/A _20386_/X VGND VGND VPWR VPWR _23410_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15025__A2_N _15024_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22128_ _21064_/X _22124_/X _22127_/X VGND VGND VPWR VPWR _22128_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_26_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14950_ _14950_/A VGND VGND VPWR VPWR _14950_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22059_ _14734_/Y _19614_/A _22060_/A _19610_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_89_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13901_ _13900_/X VGND VGND VPWR VPWR _15435_/B sky130_fd_sc_hd__buf_2
XFILLER_48_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14881_ _14873_/B _14880_/X VGND VGND VPWR VPWR _14881_/Y sky130_fd_sc_hd__nor2_4
XFILLER_208_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15065__A2 _14996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ _13564_/Y _13831_/X _11809_/X _13831_/X VGND VGND VPWR VPWR _13832_/X sky130_fd_sc_hd__a2bb2o_4
X_16620_ _16620_/A VGND VGND VPWR VPWR _16620_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16551_ _15718_/A VGND VGND VPWR VPWR _16552_/A sky130_fd_sc_hd__buf_2
XANTENNA__21481__A _21676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13763_ _25284_/Q VGND VGND VPWR VPWR _14706_/A sky130_fd_sc_hd__inv_2
XFILLER_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12823__B2 _22755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _12729_/A _12713_/X VGND VGND VPWR VPWR _12731_/A sky130_fd_sc_hd__or2_4
X_15502_ _11727_/A _15500_/X HADDR[23] _15500_/X VGND VGND VPWR VPWR _15502_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16482_ _16482_/A VGND VGND VPWR VPWR _16482_/Y sky130_fd_sc_hd__inv_2
X_19270_ _19270_/A VGND VGND VPWR VPWR _19270_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13694_ _11685_/Y _13693_/X VGND VGND VPWR VPWR _13695_/B sky130_fd_sc_hd__or2_4
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15433_ _15396_/A _15334_/D _15324_/X _15430_/Y VGND VGND VPWR VPWR _15433_/X sky130_fd_sc_hd__a211o_4
X_18221_ _18189_/A _19050_/A VGND VGND VPWR VPWR _18223_/B sky130_fd_sc_hd__or2_4
XFILLER_231_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ _12631_/C _12642_/X VGND VGND VPWR VPWR _12645_/X sky130_fd_sc_hd__or2_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15773__B1 _15636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22638__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15364_ _25002_/Q _15363_/Y VGND VGND VPWR VPWR _15364_/X sky130_fd_sc_hd__or2_4
X_18152_ _17984_/A _18152_/B VGND VGND VPWR VPWR _18152_/X sky130_fd_sc_hd__or2_4
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12576_ _25420_/Q VGND VGND VPWR VPWR _12618_/D sky130_fd_sc_hd__inv_2
XFILLER_156_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _14315_/A VGND VGND VPWR VPWR _14315_/X sky130_fd_sc_hd__buf_2
X_17103_ _17102_/X VGND VGND VPWR VPWR _17104_/B sky130_fd_sc_hd__inv_2
XFILLER_184_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18083_ _18189_/A _18083_/B VGND VGND VPWR VPWR _18083_/X sky130_fd_sc_hd__or2_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15295_ _15387_/A VGND VGND VPWR VPWR _15357_/A sky130_fd_sc_hd__inv_2
X_17034_ _17034_/A _17075_/C VGND VGND VPWR VPWR _17034_/X sky130_fd_sc_hd__or2_4
X_14246_ _14244_/Y _14245_/X _13812_/X _14245_/X VGND VGND VPWR VPWR _14246_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13439__A _13186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__B2 _21747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ _14120_/X _14176_/Y _14455_/A _14120_/X VGND VGND VPWR VPWR _25218_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12343__A _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13128_ _20776_/A _24033_/Q _20768_/A _24034_/Q VGND VGND VPWR VPWR _13128_/X sky130_fd_sc_hd__or4_4
X_18985_ _18985_/A VGND VGND VPWR VPWR _18985_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13839__B1 _11831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15654__A _15657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ _13054_/A _13053_/X _13019_/A _13055_/Y VGND VGND VPWR VPWR _13059_/X sky130_fd_sc_hd__a211o_4
X_17936_ _13550_/A _17934_/Y _17924_/B _17935_/X VGND VGND VPWR VPWR _24256_/D sky130_fd_sc_hd__o22a_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17867_ _17861_/C _17866_/X _17798_/X _17863_/B VGND VGND VPWR VPWR _17868_/A sky130_fd_sc_hd__a211o_4
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19606_ _19615_/A VGND VGND VPWR VPWR _19606_/X sky130_fd_sc_hd__buf_2
XFILLER_213_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ _24444_/Q VGND VGND VPWR VPWR _16818_/Y sky130_fd_sc_hd__inv_2
X_17798_ _16963_/Y VGND VGND VPWR VPWR _17798_/X sky130_fd_sc_hd__buf_2
XFILLER_35_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14803__A2 _13610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24851__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19537_ _21960_/B _19534_/X _11952_/X _19534_/X VGND VGND VPWR VPWR _23713_/D sky130_fd_sc_hd__a2bb2o_4
X_16749_ _15060_/Y _16748_/X _15732_/X _16748_/X VGND VGND VPWR VPWR _16749_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19468_ _18083_/B VGND VGND VPWR VPWR _19468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18950__B1 _16796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ _22312_/A _18418_/A _16261_/Y _18418_/Y VGND VGND VPWR VPWR _18419_/X sky130_fd_sc_hd__o22a_4
XFILLER_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15764__B1 _11831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19399_ _18074_/B VGND VGND VPWR VPWR _19399_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21430_ _21231_/A VGND VGND VPWR VPWR _21430_/X sky130_fd_sc_hd__buf_2
XFILLER_159_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21361_ _21361_/A _21361_/B _21358_/Y _21360_/Y VGND VGND VPWR VPWR _21361_/X sky130_fd_sc_hd__or4_4
XANTENNA__15516__B1 HADDR[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23100_ _24609_/Q _23274_/B VGND VGND VPWR VPWR _23100_/X sky130_fd_sc_hd__or2_4
X_20312_ _23439_/Q VGND VGND VPWR VPWR _20312_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24080_ _25365_/CLK _20437_/X HRESETn VGND VGND VPWR VPWR _15492_/A sky130_fd_sc_hd__dfrtp_4
X_21292_ _21060_/X _21079_/X _21292_/C _21291_/Y VGND VGND VPWR VPWR HRDATA[0] sky130_fd_sc_hd__or4_4
X_23031_ _12261_/Y _23280_/A _23030_/X VGND VGND VPWR VPWR _23031_/Y sky130_fd_sc_hd__o21ai_4
X_20243_ _11855_/A VGND VGND VPWR VPWR _20243_/X sky130_fd_sc_hd__buf_2
XFILLER_1_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20174_ _23491_/Q VGND VGND VPWR VPWR _20174_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15564__A _21172_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24982_ _24981_/CLK _15432_/X HRESETn VGND VGND VPWR VPWR _15311_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23933_ _24111_/CLK _23933_/D VGND VGND VPWR VPWR _23933_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_217_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23864_ _23577_/CLK _23864_/D VGND VGND VPWR VPWR _23864_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24592__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22815_ _22941_/A VGND VGND VPWR VPWR _22815_/X sky130_fd_sc_hd__buf_2
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23795_ _24214_/CLK _19306_/X VGND VGND VPWR VPWR _23795_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16395__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25534_ _25539_/CLK _25534_/D HRESETn VGND VGND VPWR VPWR _25534_/Q sky130_fd_sc_hd__dfrtp_4
X_22746_ _22523_/X _22744_/X _21968_/A _22745_/X VGND VGND VPWR VPWR _22746_/X sky130_fd_sc_hd__o22a_4
XFILLER_213_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18613__A1_N _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18941__B1 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25465_ _25456_/CLK _25465_/D HRESETn VGND VGND VPWR VPWR _12191_/A sky130_fd_sc_hd__dfrtp_4
X_22677_ _17257_/Y _22677_/B VGND VGND VPWR VPWR _22680_/A sky130_fd_sc_hd__or2_4
XANTENNA__12428__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12430_ _12425_/A _12425_/B _12411_/X _12427_/B VGND VGND VPWR VPWR _12430_/X sky130_fd_sc_hd__a211o_4
X_24416_ _23475_/CLK _16878_/X HRESETn VGND VGND VPWR VPWR _20108_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16953__A2_N _16952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21628_ _14761_/A _18928_/Y VGND VGND VPWR VPWR _21630_/B sky130_fd_sc_hd__or2_4
XFILLER_200_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25396_ _24812_/CLK _25396_/D HRESETn VGND VGND VPWR VPWR _12817_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12361_ _13083_/A VGND VGND VPWR VPWR _13006_/A sky130_fd_sc_hd__inv_2
X_24347_ _24354_/CLK _24347_/D HRESETn VGND VGND VPWR VPWR _24347_/Q sky130_fd_sc_hd__dfrtp_4
X_21559_ _21351_/A VGND VGND VPWR VPWR _22129_/B sky130_fd_sc_hd__buf_2
XFILLER_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14100_ _14073_/A VGND VGND VPWR VPWR _20461_/C sky130_fd_sc_hd__buf_2
XFILLER_193_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15080_ _14910_/Y _15080_/B VGND VGND VPWR VPWR _15193_/A sky130_fd_sc_hd__or2_4
X_12292_ _12218_/Y _12278_/Y _12287_/X _12291_/X VGND VGND VPWR VPWR _12292_/X sky130_fd_sc_hd__or4_4
X_24278_ _24283_/CLK _24278_/D HRESETn VGND VGND VPWR VPWR _17764_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14031_ _14042_/B VGND VGND VPWR VPWR _14031_/Y sky130_fd_sc_hd__inv_2
X_23229_ _23113_/X _23228_/X _23159_/X _24853_/Q _23115_/X VGND VGND VPWR VPWR _23229_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18770_ _18763_/A _18751_/X _18740_/X _18768_/B VGND VGND VPWR VPWR _18770_/X sky130_fd_sc_hd__a211o_4
X_15982_ _15797_/X _15977_/X _16252_/A _22608_/A _15940_/X VGND VGND VPWR VPWR _24764_/D
+ sky130_fd_sc_hd__a32o_4
X_17721_ _18289_/A _18289_/C _17720_/X VGND VGND VPWR VPWR _17721_/X sky130_fd_sc_hd__a21o_4
X_14933_ _14933_/A _14933_/B _14929_/X _14933_/D VGND VGND VPWR VPWR _14949_/C sky130_fd_sc_hd__or4_4
XANTENNA__15193__B _15294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24609__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17652_ _17641_/A _17652_/B _17652_/C VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__and3_4
XFILLER_36_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_113_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _24872_/CLK sky130_fd_sc_hd__clkbuf_1
X_14864_ _25052_/Q _14809_/B _25052_/Q _14809_/B VGND VGND VPWR VPWR _14864_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14246__B1 _13812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22308__B2 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16603_ _16603_/A VGND VGND VPWR VPWR _16603_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_176_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _25507_/CLK sky130_fd_sc_hd__clkbuf_1
X_13815_ _25277_/Q VGND VGND VPWR VPWR _13815_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14795_ _17990_/A VGND VGND VPWR VPWR _18059_/A sky130_fd_sc_hd__buf_2
X_17583_ _24299_/Q VGND VGND VPWR VPWR _17701_/A sky130_fd_sc_hd__inv_2
XANTENNA__15994__B1 _21715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19185__B1 _19184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19322_ _17958_/B VGND VGND VPWR VPWR _19322_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13746_ _25282_/Q VGND VGND VPWR VPWR _13757_/A sky130_fd_sc_hd__buf_2
X_16534_ _14423_/A VGND VGND VPWR VPWR _16534_/X sky130_fd_sc_hd__buf_2
XFILLER_232_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14549__A1 scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19253_ _23813_/Q VGND VGND VPWR VPWR _19253_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13677_ _13677_/A _13676_/X VGND VGND VPWR VPWR _20831_/B sky130_fd_sc_hd__or2_4
X_16465_ _18488_/A _16464_/X _16375_/X _16464_/X VGND VGND VPWR VPWR _24584_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15746__B1 _11797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18204_ _15703_/X _18188_/X _18203_/X _24249_/Q _18029_/A VGND VGND VPWR VPWR _18204_/X
+ sky130_fd_sc_hd__o32a_4
X_12628_ _12628_/A _12627_/X VGND VGND VPWR VPWR _12628_/X sky130_fd_sc_hd__or2_4
X_15416_ _15387_/A VGND VGND VPWR VPWR _15427_/C sky130_fd_sc_hd__buf_2
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16396_ _15099_/Y _16391_/X _16395_/X _16391_/X VGND VGND VPWR VPWR _24612_/D sky130_fd_sc_hd__a2bb2o_4
X_19184_ _19048_/A VGND VGND VPWR VPWR _19184_/X sky130_fd_sc_hd__buf_2
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15347_ _15347_/A _15346_/X VGND VGND VPWR VPWR _15352_/B sky130_fd_sc_hd__or2_4
X_18135_ _18199_/A _19200_/A VGND VGND VPWR VPWR _18135_/X sky130_fd_sc_hd__or2_4
X_12559_ _12557_/A _24869_/Q _12621_/A _12558_/Y VGND VGND VPWR VPWR _12566_/B sky130_fd_sc_hd__o22a_4
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15278_ _15259_/A _15280_/B _15277_/Y VGND VGND VPWR VPWR _15278_/X sky130_fd_sc_hd__o21a_4
X_18066_ _18168_/A _18066_/B VGND VGND VPWR VPWR _18067_/C sky130_fd_sc_hd__or2_4
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14229_ _14229_/A VGND VGND VPWR VPWR _14230_/A sky130_fd_sc_hd__buf_2
X_17017_ _16018_/Y _24404_/Q _24741_/Q _17016_/Y VGND VGND VPWR VPWR _17020_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18968_ _23913_/Q VGND VGND VPWR VPWR _18968_/Y sky130_fd_sc_hd__inv_2
X_17919_ _22005_/A VGND VGND VPWR VPWR _17919_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ _18876_/A _18890_/A _23964_/Q _24124_/Q _18893_/A VGND VGND VPWR VPWR _18899_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_226_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_72_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_72_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20930_ _20928_/Y _20924_/X _20929_/X VGND VGND VPWR VPWR _20930_/X sky130_fd_sc_hd__o21a_4
XFILLER_227_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20861_ _16713_/Y _20854_/X _20842_/X _20860_/Y VGND VGND VPWR VPWR _20861_/X sky130_fd_sc_hd__o22a_4
XFILLER_214_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15985__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22600_ _22599_/X VGND VGND VPWR VPWR _22600_/Y sky130_fd_sc_hd__inv_2
XFILLER_241_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23580_ _23475_/CLK _19927_/X VGND VGND VPWR VPWR _23580_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ _20765_/A VGND VGND VPWR VPWR _20792_/X sky130_fd_sc_hd__buf_2
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22945__A _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22531_ _15623_/Y _22531_/B VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__and2_4
XFILLER_222_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25250_ _25253_/CLK _13890_/X HRESETn VGND VGND VPWR VPWR _25250_/Q sky130_fd_sc_hd__dfrtp_4
X_22462_ _22462_/A VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__buf_2
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24201_ _24201_/CLK _24201_/D HRESETn VGND VGND VPWR VPWR _24201_/Q sky130_fd_sc_hd__dfrtp_4
X_21413_ _21409_/X _21412_/X _21251_/X VGND VGND VPWR VPWR _21413_/X sky130_fd_sc_hd__o21a_4
X_25181_ _25181_/CLK _14323_/X HRESETn VGND VGND VPWR VPWR _25181_/Q sky130_fd_sc_hd__dfrtp_4
X_22393_ _22094_/A _19923_/Y VGND VGND VPWR VPWR _22393_/X sky130_fd_sc_hd__or2_4
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14463__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24132_ _24138_/CLK _24132_/D HRESETn VGND VGND VPWR VPWR _24132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21344_ _23148_/A VGND VGND VPWR VPWR _21344_/X sky130_fd_sc_hd__buf_2
XFILLER_162_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24063_ _24431_/CLK _20909_/X HRESETn VGND VGND VPWR VPWR _24063_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17774__A _17562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21275_ _21275_/A _21275_/B _21275_/C VGND VGND VPWR VPWR _21275_/X sky130_fd_sc_hd__and3_4
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23014_ _15098_/A _23189_/B VGND VGND VPWR VPWR _23014_/X sky130_fd_sc_hd__or2_4
XFILLER_89_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20226_ _20213_/Y VGND VGND VPWR VPWR _20226_/X sky130_fd_sc_hd__buf_2
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15294__A _15294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20157_ _20155_/Y _20151_/X _20108_/X _20156_/X VGND VGND VPWR VPWR _20157_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24773__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24965_ _24339_/CLK _15468_/X HRESETn VGND VGND VPWR VPWR _13902_/A sky130_fd_sc_hd__dfrtp_4
X_20088_ _13321_/B VGND VGND VPWR VPWR _20088_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24702__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25138__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11930_ _25516_/Q _11928_/Y _11929_/Y VGND VGND VPWR VPWR _25516_/D sky130_fd_sc_hd__o21a_4
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23916_ _23916_/CLK _18962_/X VGND VGND VPWR VPWR _18958_/A sky130_fd_sc_hd__dfxtp_4
X_24896_ _24913_/CLK _15669_/X HRESETn VGND VGND VPWR VPWR _20830_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11861_ _11861_/A VGND VGND VPWR VPWR _14412_/A sky130_fd_sc_hd__buf_2
X_23847_ _24101_/CLK _23847_/D VGND VGND VPWR VPWR _19158_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_245_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14251__A1_N _14250_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23016__A _23016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_249_0_HCLK clkbuf_8_249_0_HCLK/A VGND VGND VPWR VPWR _23385_/CLK sky130_fd_sc_hd__clkbuf_1
X_13600_ _14629_/B VGND VGND VPWR VPWR _13601_/B sky130_fd_sc_hd__inv_2
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14580_/A VGND VGND VPWR VPWR _14580_/Y sky130_fd_sc_hd__inv_2
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _25544_/Q VGND VGND VPWR VPWR _11792_/Y sky130_fd_sc_hd__inv_2
X_23778_ _23850_/CLK _19354_/X VGND VGND VPWR VPWR _18055_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _14296_/A _14309_/A _25184_/Q _13531_/D VGND VGND VPWR VPWR _13532_/B sky130_fd_sc_hd__and4_4
XFILLER_186_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22729_ _22715_/X _22719_/X _22723_/X _22728_/X VGND VGND VPWR VPWR _22729_/X sky130_fd_sc_hd__or4_4
X_25517_ _23678_/CLK _25517_/D HRESETn VGND VGND VPWR VPWR _11885_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_241_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15728__B1 _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16250_ _24663_/Q VGND VGND VPWR VPWR _16250_/Y sky130_fd_sc_hd__inv_2
X_13462_ _13254_/X _13460_/X _13461_/X VGND VGND VPWR VPWR _13462_/X sky130_fd_sc_hd__and3_4
X_25448_ _25443_/CLK _12488_/Y HRESETn VGND VGND VPWR VPWR _25448_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23266__A2 _21039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15201_ _15009_/X _15078_/X _15172_/X VGND VGND VPWR VPWR _15201_/X sky130_fd_sc_hd__or3_4
X_12413_ _12412_/X VGND VGND VPWR VPWR _12413_/Y sky130_fd_sc_hd__inv_2
X_16181_ _16179_/A VGND VGND VPWR VPWR _16182_/B sky130_fd_sc_hd__buf_2
X_13393_ _13286_/X _13393_/B VGND VGND VPWR VPWR _13393_/X sky130_fd_sc_hd__or2_4
X_25379_ _25402_/CLK _25379_/D HRESETn VGND VGND VPWR VPWR _12842_/A sky130_fd_sc_hd__dfrtp_4
X_15132_ _24986_/Q VGND VGND VPWR VPWR _15399_/A sky130_fd_sc_hd__inv_2
X_12344_ _12342_/A _24827_/Q _12342_/Y _12343_/Y VGND VGND VPWR VPWR _12344_/X sky130_fd_sc_hd__o22a_4
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15063_ _15057_/X _15058_/X _15059_/X _15063_/D VGND VGND VPWR VPWR _15063_/X sky130_fd_sc_hd__or4_4
X_19940_ _19940_/A VGND VGND VPWR VPWR _19940_/Y sky130_fd_sc_hd__inv_2
X_12275_ _25468_/Q VGND VGND VPWR VPWR _12275_/Y sky130_fd_sc_hd__inv_2
X_14014_ _14014_/A VGND VGND VPWR VPWR _14015_/D sky130_fd_sc_hd__inv_2
X_19871_ _23600_/Q VGND VGND VPWR VPWR _21782_/B sky130_fd_sc_hd__inv_2
X_18822_ _18689_/A _18825_/B _18714_/X VGND VGND VPWR VPWR _18822_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_110_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18753_ _18696_/D _18753_/B VGND VGND VPWR VPWR _18756_/B sky130_fd_sc_hd__or2_4
X_15965_ HWDATA[20] VGND VGND VPWR VPWR _15965_/X sky130_fd_sc_hd__buf_2
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17704_ _17701_/B _17704_/B _17702_/C VGND VGND VPWR VPWR _17704_/X sky130_fd_sc_hd__and3_4
Xclkbuf_6_59_0_HCLK clkbuf_6_58_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14916_ _25013_/Q VGND VGND VPWR VPWR _14916_/Y sky130_fd_sc_hd__inv_2
X_18684_ _18604_/A VGND VGND VPWR VPWR _18797_/A sky130_fd_sc_hd__inv_2
X_15896_ _15896_/A VGND VGND VPWR VPWR _15896_/X sky130_fd_sc_hd__buf_2
XFILLER_36_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _17567_/Y _17590_/X VGND VGND VPWR VPWR _17635_/X sky130_fd_sc_hd__or2_4
X_14847_ _14811_/C _14825_/X _14811_/C _14825_/X VGND VGND VPWR VPWR _14848_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13452__A _13420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17566_ _24326_/Q VGND VGND VPWR VPWR _17566_/Y sky130_fd_sc_hd__inv_2
X_14778_ _13597_/X VGND VGND VPWR VPWR _14778_/X sky130_fd_sc_hd__buf_2
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14267__B _14232_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15982__A3 _16252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19305_ _19148_/A VGND VGND VPWR VPWR _19305_/X sky130_fd_sc_hd__buf_2
X_16517_ _16517_/A VGND VGND VPWR VPWR _16517_/Y sky130_fd_sc_hd__inv_2
X_13729_ _11672_/Y _13695_/B VGND VGND VPWR VPWR _13729_/Y sky130_fd_sc_hd__nand2_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17497_ _17496_/X VGND VGND VPWR VPWR _17497_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19236_ _19249_/A VGND VGND VPWR VPWR _19236_/X sky130_fd_sc_hd__buf_2
XFILLER_231_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16448_ _24588_/Q VGND VGND VPWR VPWR _16448_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16392__B1 _16389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17578__B _17578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19167_ _19166_/X VGND VGND VPWR VPWR _19181_/A sky130_fd_sc_hd__inv_2
XANTENNA__16913__D _16912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16379_ _16379_/A VGND VGND VPWR VPWR _22459_/A sky130_fd_sc_hd__buf_2
XANTENNA__25231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18118_ _17979_/A _18118_/B VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__or2_4
XANTENNA__16144__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19098_ _13774_/X _13775_/X _13744_/X _20149_/B VGND VGND VPWR VPWR _19099_/A sky130_fd_sc_hd__or4_4
XFILLER_172_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18049_ _18234_/A _18045_/X _18049_/C VGND VGND VPWR VPWR _18049_/X sky130_fd_sc_hd__or3_4
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21060_ _21060_/A _21060_/B _21060_/C VGND VGND VPWR VPWR _21060_/X sky130_fd_sc_hd__and3_4
XFILLER_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20011_ _21497_/B _20006_/X _20010_/X _20006_/X VGND VGND VPWR VPWR _20011_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16447__B2 _16446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16003__A _16003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16970__A1_N _24727_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24750_ _24738_/CLK _16013_/X HRESETn VGND VGND VPWR VPWR _16010_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_239_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21962_ _21941_/A _21962_/B VGND VGND VPWR VPWR _21962_/X sky130_fd_sc_hd__or2_4
XANTENNA__24113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _23669_/CLK _23701_/D VGND VGND VPWR VPWR _23701_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16355__A1_N _16354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20913_ _20900_/X _20912_/Y _24501_/Q _20904_/X VGND VGND VPWR VPWR _20913_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24681_ _24657_/CLK _16204_/X HRESETn VGND VGND VPWR VPWR _16201_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15958__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21893_ _21893_/A _21892_/X VGND VGND VPWR VPWR _21893_/X sky130_fd_sc_hd__and2_4
XFILLER_227_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23615_/CLK _23632_/D VGND VGND VPWR VPWR _13371_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _16723_/Y _20833_/X _20842_/X _20843_/X VGND VGND VPWR VPWR _20845_/A sky130_fd_sc_hd__o22a_4
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_16_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _23678_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _23563_/CLK _19970_/X VGND VGND VPWR VPWR _23563_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17769__A _17762_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20775_ _24033_/Q VGND VGND VPWR VPWR _20775_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25302_ _24196_/CLK _13684_/X HRESETn VGND VGND VPWR VPWR _25302_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_79_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24757_/CLK sky130_fd_sc_hd__clkbuf_1
X_22514_ _16608_/Y _22460_/X _21591_/X _22513_/X VGND VGND VPWR VPWR _22514_/X sky130_fd_sc_hd__o22a_4
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _23494_/CLK _20166_/X VGND VGND VPWR VPWR _23494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25233_ _25105_/CLK _25233_/D HRESETn VGND VGND VPWR VPWR _13994_/B sky130_fd_sc_hd__dfrtp_4
X_22445_ _16156_/Y _22444_/X _22440_/X _11837_/Y _22283_/X VGND VGND VPWR VPWR _22445_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_155_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22456__B1 _25446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19321__B1 _19254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25164_ _24121_/CLK _14372_/X HRESETn VGND VGND VPWR VPWR _25164_/Q sky130_fd_sc_hd__dfrtp_4
X_22376_ _22380_/A _22374_/X _22376_/C VGND VGND VPWR VPWR _22376_/X sky130_fd_sc_hd__and3_4
XFILLER_135_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24115_ _25145_/CLK _20980_/X HRESETn VGND VGND VPWR VPWR _24115_/Q sky130_fd_sc_hd__dfrtp_4
X_21327_ _16731_/Y VGND VGND VPWR VPWR _22171_/A sky130_fd_sc_hd__buf_2
X_25095_ _25093_/CLK _25095_/D HRESETn VGND VGND VPWR VPWR _14568_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22759__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ _15791_/C VGND VGND VPWR VPWR _16190_/C sky130_fd_sc_hd__buf_2
X_24046_ _24915_/CLK _20829_/X HRESETn VGND VGND VPWR VPWR _13147_/A sky130_fd_sc_hd__dfrtp_4
X_21258_ _21248_/A VGND VGND VPWR VPWR _21259_/A sky130_fd_sc_hd__buf_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20209_ _23477_/Q VGND VGND VPWR VPWR _20209_/Y sky130_fd_sc_hd__inv_2
X_21189_ _21183_/X _21188_/X _17729_/Y VGND VGND VPWR VPWR _21189_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14449__B1 _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19388__B1 _19254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15752__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12962_ _12961_/X VGND VGND VPWR VPWR _12962_/Y sky130_fd_sc_hd__inv_2
X_15750_ _15737_/X _15722_/X _15748_/X _24876_/Q _15749_/X VGND VGND VPWR VPWR _24876_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_246_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24948_ _23407_/CLK _15511_/X HRESETn VGND VGND VPWR VPWR _11736_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_218_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11913_ _11913_/A VGND VGND VPWR VPWR _11913_/Y sky130_fd_sc_hd__inv_2
X_14701_ _14700_/X VGND VGND VPWR VPWR _22228_/A sky130_fd_sc_hd__buf_2
XANTENNA__15471__B _14232_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12893_ _12891_/X _12888_/B _12893_/C VGND VGND VPWR VPWR _12894_/A sky130_fd_sc_hd__or3_4
X_15681_ _22738_/A VGND VGND VPWR VPWR _15681_/X sky130_fd_sc_hd__buf_2
XANTENNA__15949__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24879_ _24889_/CLK _15745_/X HRESETn VGND VGND VPWR VPWR _24879_/Q sky130_fd_sc_hd__dfrtp_4
X_17420_ _24086_/Q _13976_/Y _21018_/A _13976_/A VGND VGND VPWR VPWR _17420_/X sky130_fd_sc_hd__o22a_4
X_11844_ _25531_/Q VGND VGND VPWR VPWR _11844_/Y sky130_fd_sc_hd__inv_2
X_14632_ _14639_/A _14639_/B _14631_/Y VGND VGND VPWR VPWR _14632_/X sky130_fd_sc_hd__a21o_4
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _25103_/Q VGND VGND VPWR VPWR _14563_/Y sky130_fd_sc_hd__inv_2
X_17351_ _17258_/Y _17345_/X _17298_/A _17348_/B VGND VGND VPWR VPWR _17351_/X sky130_fd_sc_hd__a211o_4
XFILLER_214_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _25549_/Q VGND VGND VPWR VPWR _11775_/Y sky130_fd_sc_hd__inv_2
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _24644_/Q VGND VGND VPWR VPWR _16302_/Y sky130_fd_sc_hd__inv_2
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _13514_/A VGND VGND VPWR VPWR _13514_/Y sky130_fd_sc_hd__inv_2
X_14494_ _14494_/A VGND VGND VPWR VPWR _21726_/A sky130_fd_sc_hd__inv_2
X_17282_ _17282_/A VGND VGND VPWR VPWR _24376_/D sky130_fd_sc_hd__inv_2
XFILLER_186_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19021_ _19019_/Y _19020_/X _18975_/X _19020_/X VGND VGND VPWR VPWR _23895_/D sky130_fd_sc_hd__a2bb2o_4
X_13445_ _13413_/A _23813_/Q VGND VGND VPWR VPWR _13445_/X sky130_fd_sc_hd__or2_4
X_16233_ _24668_/Q VGND VGND VPWR VPWR _16233_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15199__A _14996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19312__B1 _19220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13376_ _13209_/X _13360_/X _13375_/X _25335_/Q _11974_/X VGND VGND VPWR VPWR _13376_/X
+ sky130_fd_sc_hd__o32a_4
X_16164_ _22162_/A VGND VGND VPWR VPWR _16164_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16126__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20833__A _20854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12327_ _12327_/A VGND VGND VPWR VPWR _12327_/Y sky130_fd_sc_hd__inv_2
X_15115_ _24988_/Q _15114_/A _15401_/A _15114_/Y VGND VGND VPWR VPWR _15116_/D sky130_fd_sc_hd__o22a_4
X_16095_ _11730_/Y _22513_/B VGND VGND VPWR VPWR _16096_/A sky130_fd_sc_hd__and2_4
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24695__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15046_ _15259_/A _24458_/Q _15259_/A _24458_/Q VGND VGND VPWR VPWR _15049_/C sky130_fd_sc_hd__a2bb2o_4
X_19923_ _23580_/Q VGND VGND VPWR VPWR _19923_/Y sky130_fd_sc_hd__inv_2
X_12258_ _12294_/A VGND VGND VPWR VPWR _12464_/A sky130_fd_sc_hd__buf_2
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24624__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19854_ _19853_/Y _19851_/X _19810_/X _19851_/X VGND VGND VPWR VPWR _19854_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12189_ _12397_/A _24784_/Q _12397_/A _24784_/Q VGND VGND VPWR VPWR _12189_/X sky130_fd_sc_hd__a2bb2o_4
X_18805_ _18805_/A _18805_/B VGND VGND VPWR VPWR _18805_/X sky130_fd_sc_hd__or2_4
X_19785_ _19784_/Y _19780_/X _19761_/X _19765_/Y VGND VGND VPWR VPWR _19785_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17861__B _17861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16997_ _24739_/Q _16996_/A _16038_/Y _16996_/Y VGND VGND VPWR VPWR _16998_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16758__A _16762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15662__A _15661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18736_ _18736_/A VGND VGND VPWR VPWR _18736_/Y sky130_fd_sc_hd__inv_2
X_15948_ HWDATA[29] VGND VGND VPWR VPWR _15948_/X sky130_fd_sc_hd__buf_2
XFILLER_110_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18667_ _18660_/X _18662_/X _18664_/X _18666_/X VGND VGND VPWR VPWR _18667_/X sky130_fd_sc_hd__or4_4
X_15879_ _12829_/Y _15877_/X _11763_/X _15877_/X VGND VGND VPWR VPWR _24818_/D sky130_fd_sc_hd__a2bb2o_4
X_17618_ _17610_/B _17610_/D _17610_/A VGND VGND VPWR VPWR _17618_/X sky130_fd_sc_hd__o21a_4
X_18598_ _18598_/A _18597_/Y _18598_/C VGND VGND VPWR VPWR _18598_/X sky130_fd_sc_hd__and3_4
XANTENNA__25483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22495__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15955__A3 HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_232_0_HCLK clkbuf_7_116_0_HCLK/X VGND VGND VPWR VPWR _23970_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14711__A1_N _14709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17549_ _24324_/Q VGND VGND VPWR VPWR _17569_/A sky130_fd_sc_hd__inv_2
XFILLER_149_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20560_ _23951_/Q _18877_/X VGND VGND VPWR VPWR _20561_/B sky130_fd_sc_hd__nand2_4
XANTENNA__23103__B _23100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20161__B2 _20156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19219_ _18104_/B VGND VGND VPWR VPWR _19219_/Y sky130_fd_sc_hd__inv_2
X_20491_ _20490_/X VGND VGND VPWR VPWR _23976_/D sky130_fd_sc_hd__buf_2
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22230_ _22226_/A _22230_/B VGND VGND VPWR VPWR _22230_/X sky130_fd_sc_hd__or2_4
XFILLER_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16117__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21839__A _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14391__A2 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21110__B1 _21882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19854__B2 _19851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22661__C _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22161_ _21449_/A _22160_/X VGND VGND VPWR VPWR _22161_/X sky130_fd_sc_hd__and2_4
XFILLER_161_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21112_ _24721_/Q _21067_/X _21101_/X _21111_/X VGND VGND VPWR VPWR _21112_/X sky130_fd_sc_hd__a211o_4
XFILLER_105_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22092_ _22087_/X _22091_/X _14686_/X VGND VGND VPWR VPWR _22092_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_114_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21043_ _21043_/A VGND VGND VPWR VPWR _21058_/A sky130_fd_sc_hd__buf_2
XFILLER_247_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21574__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17771__B _16952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25472__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24802_ _24794_/CLK _15901_/X HRESETn VGND VGND VPWR VPWR _22641_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15572__A _15584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22994_ _22994_/A _22882_/X VGND VGND VPWR VPWR _22994_/X sky130_fd_sc_hd__or2_4
XFILLER_228_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21945_ _21945_/A _21945_/B _21945_/C VGND VGND VPWR VPWR _21945_/X sky130_fd_sc_hd__and3_4
X_24733_ _24735_/CLK _24733_/D HRESETn VGND VGND VPWR VPWR _16053_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13804__B _16464_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24100__D _20970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24657_/CLK _24664_/D HRESETn VGND VGND VPWR VPWR _24664_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_203_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _21235_/X VGND VGND VPWR VPWR _22299_/B sky130_fd_sc_hd__buf_2
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23615_/CLK _19830_/X VGND VGND VPWR VPWR _23615_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20825_/Y _20826_/Y _13147_/B VGND VGND VPWR VPWR _20827_/X sky130_fd_sc_hd__o21a_4
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ _24592_/CLK _24595_/D HRESETn VGND VGND VPWR VPWR _15095_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18345__A1 _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23546_ _23684_/CLK _20023_/X VGND VGND VPWR VPWR _20021_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20758_ _13142_/D _20753_/X VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__or2_4
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _23400_/CLK _23477_/D VGND VGND VPWR VPWR _23477_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20689_ _20499_/X _20506_/X _20621_/B VGND VGND VPWR VPWR _24008_/D sky130_fd_sc_hd__o21a_4
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16862__A1_N _14946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13271_/A VGND VGND VPWR VPWR _13317_/A sky130_fd_sc_hd__buf_2
X_25216_ _25215_/CLK _25216_/D HRESETn VGND VGND VPWR VPWR _14174_/B sky130_fd_sc_hd__dfrtp_4
X_22428_ _22428_/A _21091_/B VGND VGND VPWR VPWR _22428_/X sky130_fd_sc_hd__or2_4
XANTENNA__19845__B2 _19844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13161_ _13443_/A VGND VGND VPWR VPWR _13192_/A sky130_fd_sc_hd__buf_2
X_25147_ _25223_/CLK _14431_/X HRESETn VGND VGND VPWR VPWR _14430_/A sky130_fd_sc_hd__dfstp_4
X_22359_ _21945_/A _22357_/X _22358_/X VGND VGND VPWR VPWR _22359_/X sky130_fd_sc_hd__and3_4
XFILLER_109_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18123__A _18234_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12112_ _12101_/Y _12111_/X _11834_/X _12111_/X VGND VGND VPWR VPWR _25483_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13092_ _12386_/Y _13107_/B VGND VGND VPWR VPWR _13092_/X sky130_fd_sc_hd__or2_4
X_25078_ _23836_/CLK _25078_/D HRESETn VGND VGND VPWR VPWR _13611_/A sky130_fd_sc_hd__dfrtp_4
X_12043_ _12050_/A VGND VGND VPWR VPWR _12043_/X sky130_fd_sc_hd__buf_2
X_16920_ _24270_/Q VGND VGND VPWR VPWR _16920_/Y sky130_fd_sc_hd__inv_2
X_24029_ _24029_/CLK _24029_/D HRESETn VGND VGND VPWR VPWR _13142_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12171__A _14342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_249_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21484__A _21676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16851_ _14925_/Y _16849_/X _16613_/X _16849_/X VGND VGND VPWR VPWR _24427_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16578__A _16578_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22299__B _22299_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15802_ _15802_/A VGND VGND VPWR VPWR _15802_/X sky130_fd_sc_hd__buf_2
X_19570_ _23701_/Q VGND VGND VPWR VPWR _19570_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16782_ _16782_/A VGND VGND VPWR VPWR _16782_/X sky130_fd_sc_hd__buf_2
X_13994_ _13994_/A _13994_/B VGND VGND VPWR VPWR _14032_/B sky130_fd_sc_hd__or2_4
XFILLER_207_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18521_ _18492_/A _18517_/X _18521_/C VGND VGND VPWR VPWR _18521_/X sky130_fd_sc_hd__and3_4
X_15733_ _15557_/X _15722_/X _15732_/X _24886_/Q _15720_/X VGND VGND VPWR VPWR _24886_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12945_ _12927_/A _12943_/X _12945_/C VGND VGND VPWR VPWR _25386_/D sky130_fd_sc_hd__and3_4
XFILLER_218_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19781__B1 _19734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18452_ _16271_/Y _24166_/Q _21340_/A _18433_/Y VGND VGND VPWR VPWR _18452_/X sky130_fd_sc_hd__a2bb2o_4
X_15664_ _15663_/X VGND VGND VPWR VPWR _15664_/X sky130_fd_sc_hd__buf_2
XANTENNA__16595__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _12839_/Y _12873_/X _12868_/B _12875_/X VGND VGND VPWR VPWR _12876_/X sky130_fd_sc_hd__a211o_4
XFILLER_34_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15937__A3 _15933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _23994_/Q _20653_/A VGND VGND VPWR VPWR _17404_/B sky130_fd_sc_hd__or2_4
XFILLER_233_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _13582_/Y _14571_/B VGND VGND VPWR VPWR _14615_/Y sky130_fd_sc_hd__nand2_4
X_11827_ _16252_/A VGND VGND VPWR VPWR _11827_/X sky130_fd_sc_hd__buf_2
X_18383_ _24201_/Q VGND VGND VPWR VPWR _18383_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _23003_/A _15590_/X _11787_/X _15590_/X VGND VGND VPWR VPWR _15595_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17212_/A _17333_/Y VGND VGND VPWR VPWR _17334_/X sky130_fd_sc_hd__or2_4
XFILLER_159_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ HWDATA[29] VGND VGND VPWR VPWR _11758_/X sky130_fd_sc_hd__buf_2
X_14546_ _13993_/X _14545_/Y _14004_/X VGND VGND VPWR VPWR _14546_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16347__B1 _16252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_62_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _25103_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _17256_/X _17265_/B VGND VGND VPWR VPWR _17265_/X sky130_fd_sc_hd__or2_4
XANTENNA__16898__B2 _14791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11689_ _24241_/Q VGND VGND VPWR VPWR _22550_/A sky130_fd_sc_hd__inv_2
X_14477_ _25128_/Q VGND VGND VPWR VPWR _14477_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21891__B2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12346__A _24843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19004_ _19020_/A VGND VGND VPWR VPWR _19004_/X sky130_fd_sc_hd__buf_2
XANTENNA__24876__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16216_ _16214_/Y _16210_/X _15957_/X _16215_/X VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__a2bb2o_4
X_13428_ _13428_/A _13428_/B VGND VGND VPWR VPWR _13430_/B sky130_fd_sc_hd__or2_4
X_17196_ _23091_/A _17195_/A _16311_/Y _17248_/B VGND VGND VPWR VPWR _17196_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18639__A2 _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24805__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24962__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12384__B2 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13359_ _13391_/A _13359_/B _13359_/C VGND VGND VPWR VPWR _13360_/C sky130_fd_sc_hd__or3_4
X_16147_ _22613_/A VGND VGND VPWR VPWR _16147_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22840__B1 _17832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15657__A _15657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16078_ _16078_/A VGND VGND VPWR VPWR _16078_/Y sky130_fd_sc_hd__inv_2
X_15029_ _15250_/A _24464_/Q _15251_/A _22682_/A VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__o22a_4
X_19906_ _19902_/Y _19905_/X _19626_/X _19905_/X VGND VGND VPWR VPWR _23588_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12081__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19837_ _19837_/A _13771_/X _18914_/X VGND VGND VPWR VPWR _19838_/A sky130_fd_sc_hd__or3_4
XANTENNA__16488__A _16495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19768_ _13260_/B VGND VGND VPWR VPWR _19768_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21159__B1 _14890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22002__B _21880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18719_ _24160_/Q _18719_/B VGND VGND VPWR VPWR _18719_/X sky130_fd_sc_hd__or2_4
Xclkbuf_5_29_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ _19698_/Y VGND VGND VPWR VPWR _19699_/X sky130_fd_sc_hd__buf_2
X_21730_ _21730_/A _21730_/B _21730_/C _21729_/X VGND VGND VPWR VPWR _21731_/B sky130_fd_sc_hd__and4_4
XFILLER_25_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21841__B _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21661_ _13748_/A _21660_/X VGND VGND VPWR VPWR _21661_/Y sky130_fd_sc_hd__nor2_4
X_23400_ _23400_/CLK _23400_/D VGND VGND VPWR VPWR _20413_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_212_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18208__A _18102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23320__A1 _21547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20612_ _20448_/X VGND VGND VPWR VPWR _20612_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23320__B2 _22851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24380_ _24383_/CLK _17169_/X HRESETn VGND VGND VPWR VPWR _24380_/Q sky130_fd_sc_hd__dfrtp_4
X_21592_ _21592_/A VGND VGND VPWR VPWR _21752_/B sky130_fd_sc_hd__buf_2
XFILLER_178_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22674__A3 _22148_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23331_ _23299_/A _23331_/B _23331_/C _23330_/X VGND VGND VPWR VPWR _23331_/X sky130_fd_sc_hd__or4_4
X_20543_ _24085_/Q _20543_/B VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__and2_4
XFILLER_20_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23262_ _16558_/A _22411_/X _15676_/X _23261_/X VGND VGND VPWR VPWR _23263_/C sky130_fd_sc_hd__a211o_4
X_20474_ _20445_/A _20442_/A VGND VGND VPWR VPWR _20477_/C sky130_fd_sc_hd__and2_4
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17766__B _17766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25001_ _25002_/CLK _25001_/D HRESETn VGND VGND VPWR VPWR _25001_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22213_ _21260_/A _22213_/B _22212_/X VGND VGND VPWR VPWR _22214_/C sky130_fd_sc_hd__and3_4
XFILLER_192_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23193_ _23188_/X _23189_/X _23192_/X VGND VGND VPWR VPWR _23194_/D sky130_fd_sc_hd__and3_4
XFILLER_134_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22144_ _22144_/A VGND VGND VPWR VPWR _22145_/C sky130_fd_sc_hd__buf_2
XFILLER_105_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17782__A _16925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22075_ _22380_/A _22072_/X _22075_/C VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__and3_4
XFILLER_126_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13875__A1 _20681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21026_ _25304_/Q _21026_/B VGND VGND VPWR VPWR _21026_/X sky130_fd_sc_hd__and2_4
XFILLER_48_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12313__A2_N _24841_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22977_ _22976_/X VGND VGND VPWR VPWR _22977_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22898__B1 _22816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12730_ _12730_/A VGND VGND VPWR VPWR _12741_/C sky130_fd_sc_hd__buf_2
X_24716_ _24689_/CLK _16101_/X HRESETn VGND VGND VPWR VPWR _23296_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21928_ _22237_/A _21920_/X _21927_/X VGND VGND VPWR VPWR _21928_/X sky130_fd_sc_hd__or3_4
XANTENNA__16577__B1 _16407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18030__A3 _18028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12661_ _12616_/B _12669_/B VGND VGND VPWR VPWR _12666_/B sky130_fd_sc_hd__or2_4
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _25111_/Q _22129_/B VGND VGND VPWR VPWR _21863_/B sky130_fd_sc_hd__nand2_4
X_24647_ _24641_/CLK _24647_/D HRESETn VGND VGND VPWR VPWR _24647_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14400_/A VGND VGND VPWR VPWR _14400_/X sky130_fd_sc_hd__buf_2
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12590_/Y _24864_/Q _25434_/Q _12591_/Y VGND VGND VPWR VPWR _12598_/B sky130_fd_sc_hd__a2bb2o_4
X_15380_ _15380_/A _15384_/B VGND VGND VPWR VPWR _15380_/Y sky130_fd_sc_hd__nand2_4
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24578_ _24562_/CLK _16484_/X HRESETn VGND VGND VPWR VPWR _16482_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _14315_/A _14330_/X _25323_/Q _14320_/A VGND VGND VPWR VPWR _14331_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_49_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_49_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _23529_/CLK _20068_/X VGND VGND VPWR VPWR _20067_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11810__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16861__A _19091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14256_/Y _14261_/Y sda_oen_o_S5 _14256_/Y VGND VGND VPWR VPWR _14262_/X
+ sky130_fd_sc_hd__a2bb2o_4
X_17050_ _17048_/Y _17137_/B _17050_/C _17050_/D VGND VGND VPWR VPWR _17054_/B sky130_fd_sc_hd__or4_4
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15552__B2 _15547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22417__A3 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _13417_/A _13213_/B VGND VGND VPWR VPWR _13213_/X sky130_fd_sc_hd__or2_4
X_16001_ _14199_/A _16000_/X VGND VGND VPWR VPWR _16001_/X sky130_fd_sc_hd__or2_4
XANTENNA__17829__B1 _16964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14193_ _14192_/X VGND VGND VPWR VPWR _14193_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13144_ _13143_/X VGND VGND VPWR VPWR _13144_/X sky130_fd_sc_hd__buf_2
XFILLER_152_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16501__B1 _16414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15855__A2 _15774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13075_ _12367_/A _13074_/Y VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__or2_4
X_17952_ _17941_/A _17950_/X _17952_/C VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__and3_4
XFILLER_183_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12026_ _24108_/Q _12003_/X _12025_/Y VGND VGND VPWR VPWR _20976_/A sky130_fd_sc_hd__o21a_4
X_16903_ _16113_/Y _17752_/A _16113_/Y _17752_/A VGND VGND VPWR VPWR _16904_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11877__B1 _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18254__B1 _11830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17883_ _16937_/A _17883_/B VGND VGND VPWR VPWR _17883_/X sky130_fd_sc_hd__or2_4
X_19622_ _23684_/Q VGND VGND VPWR VPWR _19622_/Y sky130_fd_sc_hd__inv_2
X_16834_ _16853_/A VGND VGND VPWR VPWR _16834_/X sky130_fd_sc_hd__buf_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19553_ _19547_/Y _19552_/X _19439_/X _19552_/X VGND VGND VPWR VPWR _23708_/D sky130_fd_sc_hd__a2bb2o_4
X_16765_ _16764_/Y _16762_/X _16417_/X _16762_/X VGND VGND VPWR VPWR _16765_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13977_ _13962_/X VGND VGND VPWR VPWR _13977_/Y sky130_fd_sc_hd__inv_2
X_18504_ _18487_/A _18486_/X _18510_/A _18503_/X VGND VGND VPWR VPWR _18504_/X sky130_fd_sc_hd__or4_4
XANTENNA__19754__B1 _19753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15716_ _15715_/X VGND VGND VPWR VPWR _22146_/B sky130_fd_sc_hd__buf_2
X_12928_ _12924_/X VGND VGND VPWR VPWR _12929_/B sky130_fd_sc_hd__inv_2
X_19484_ _19483_/Y VGND VGND VPWR VPWR _19484_/X sky130_fd_sc_hd__buf_2
XANTENNA__16568__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21661__B _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16696_ _16696_/A VGND VGND VPWR VPWR _16696_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21561__B1 _14178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18435_ _21340_/A _18433_/Y _22107_/A _18482_/A VGND VGND VPWR VPWR _18435_/X sky130_fd_sc_hd__a2bb2o_4
X_15647_ _15647_/A VGND VGND VPWR VPWR _15647_/Y sky130_fd_sc_hd__inv_2
X_12859_ _12773_/Y _12819_/Y _12787_/Y _12762_/A VGND VGND VPWR VPWR _12859_/X sky130_fd_sc_hd__or4_4
XANTENNA__18309__A1 _18306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18028__A _18069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16139__A1_N _16138_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18366_ _18366_/A VGND VGND VPWR VPWR _18366_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15578_ _23245_/A _15572_/X _11763_/X _15577_/X VGND VGND VPWR VPWR _15578_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20116__B2 _20109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17317_ _17341_/A _17338_/A _17317_/C VGND VGND VPWR VPWR _17326_/D sky130_fd_sc_hd__or3_4
X_14529_ _14524_/A _14528_/X _14487_/A _14526_/X VGND VGND VPWR VPWR _14529_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11801__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18297_ _21834_/A _18288_/X _17710_/X VGND VGND VPWR VPWR _18297_/X sky130_fd_sc_hd__a21o_4
XFILLER_175_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ _17305_/A _17248_/B VGND VGND VPWR VPWR _17248_/X sky130_fd_sc_hd__or2_4
XANTENNA__23066__B1 _17751_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16740__B1 _16385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15543__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12357__B2 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20294__A2_N _20291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_6_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _24623_/Q _17378_/A _16302_/Y _17293_/A VGND VGND VPWR VPWR _17179_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_227_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20190_ _20190_/A VGND VGND VPWR VPWR _20190_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15846__A2 _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11868__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22900_ _22944_/A _22900_/B _22900_/C VGND VGND VPWR VPWR _22900_/X sky130_fd_sc_hd__and3_4
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23880_ _23880_/CLK _23880_/D VGND VGND VPWR VPWR _19065_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_229_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22831_ _24537_/Q _22541_/X _22542_/X _22830_/X VGND VGND VPWR VPWR _22831_/X sky130_fd_sc_hd__a211o_4
XFILLER_244_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22762_ _21082_/A _22759_/X _22723_/A _22761_/X VGND VGND VPWR VPWR _22762_/Y sky130_fd_sc_hd__a22oi_4
X_25550_ _24697_/CLK _11774_/X HRESETn VGND VGND VPWR VPWR _25550_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21713_ _21530_/X _21712_/X _21532_/X _24863_/Q _21538_/X VGND VGND VPWR VPWR _21714_/B
+ sky130_fd_sc_hd__a32o_4
X_24501_ _24532_/CLK _16688_/X HRESETn VGND VGND VPWR VPWR _24501_/Q sky130_fd_sc_hd__dfrtp_4
X_25481_ _24196_/CLK _12117_/X HRESETn VGND VGND VPWR VPWR _25481_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _22692_/X VGND VGND VPWR VPWR _22693_/Y sky130_fd_sc_hd__inv_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24798__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21644_ _21644_/A _21644_/B VGND VGND VPWR VPWR _21644_/X sky130_fd_sc_hd__or2_4
X_24432_ _24431_/CLK _16842_/X HRESETn VGND VGND VPWR VPWR _16841_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24727__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24363_ _24346_/CLK _24363_/D HRESETn VGND VGND VPWR VPWR _17212_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17777__A _23332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _16273_/Y _16192_/A _15124_/A _16731_/Y VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__a2bb2o_4
X_23314_ _15026_/A _22673_/B _23190_/X VGND VGND VPWR VPWR _23314_/X sky130_fd_sc_hd__o21a_4
X_20526_ _20524_/X _20525_/X _20620_/A VGND VGND VPWR VPWR _20526_/X sky130_fd_sc_hd__o21a_4
X_24294_ _24272_/CLK _17779_/X HRESETn VGND VGND VPWR VPWR _23332_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_181_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15534__B2 _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23245_ _23245_/A _22890_/B VGND VGND VPWR VPWR _23245_/X sky130_fd_sc_hd__and2_4
XANTENNA__15297__A _15293_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20457_ _23940_/Q VGND VGND VPWR VPWR _20457_/X sky130_fd_sc_hd__buf_2
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22280__A1 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23176_ _23174_/X _23176_/B _22929_/X VGND VGND VPWR VPWR _23176_/X sky130_fd_sc_hd__or3_4
X_20388_ _20388_/A VGND VGND VPWR VPWR _22252_/B sky130_fd_sc_hd__inv_2
XFILLER_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22127_ _21578_/X _22125_/X _21584_/X _22126_/X VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22058_ _22058_/A VGND VGND VPWR VPWR _22058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13900_ _13942_/A _13934_/A _13899_/X VGND VGND VPWR VPWR _13900_/X sky130_fd_sc_hd__or3_4
X_21009_ _21008_/A _21008_/B _24341_/Q _21008_/X VGND VGND VPWR VPWR _23983_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12520__B2 _24871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14880_ _14879_/X VGND VGND VPWR VPWR _14880_/X sky130_fd_sc_hd__buf_2
XANTENNA__16798__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18251__A3 _16248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22858__A _21881_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21762__A _21731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _13838_/A VGND VGND VPWR VPWR _13831_/X sky130_fd_sc_hd__buf_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16856__A _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12267__A2_N _24779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16550_ _16550_/A VGND VGND VPWR VPWR _16550_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13762_ _25285_/Q VGND VGND VPWR VPWR _13762_/X sky130_fd_sc_hd__buf_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_204_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15501_ _11718_/A _15500_/X HWRITE _15500_/X VGND VGND VPWR VPWR _24954_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12713_ _12713_/A _12732_/A VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__or2_4
X_16481_ _16480_/Y _16476_/X _16395_/X _16476_/X VGND VGND VPWR VPWR _24579_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_243_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13693_ _13693_/A _13692_/X VGND VGND VPWR VPWR _13693_/X sky130_fd_sc_hd__or2_4
XFILLER_188_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18220_ _13639_/X _18220_/B _18220_/C VGND VGND VPWR VPWR _18220_/X sky130_fd_sc_hd__and3_4
X_15432_ _15424_/B _15432_/B _15427_/C VGND VGND VPWR VPWR _15432_/X sky130_fd_sc_hd__and3_4
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12644_ _12644_/A _12644_/B VGND VGND VPWR VPWR _12646_/B sky130_fd_sc_hd__or2_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18790__B _18733_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18151_ _14656_/A _18149_/X _18150_/X VGND VGND VPWR VPWR _18151_/X sky130_fd_sc_hd__and3_4
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _12574_/Y _24872_/Q _12574_/Y _24872_/Q VGND VGND VPWR VPWR _12578_/C sky130_fd_sc_hd__a2bb2o_4
X_15363_ _15363_/A VGND VGND VPWR VPWR _15363_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21846__B2 _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _17016_/Y _17101_/X VGND VGND VPWR VPWR _17102_/X sky130_fd_sc_hd__or2_4
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _14320_/A VGND VGND VPWR VPWR _14315_/A sky130_fd_sc_hd__inv_2
X_18082_ _17991_/X _18082_/B _18082_/C VGND VGND VPWR VPWR _18082_/X sky130_fd_sc_hd__and3_4
XFILLER_172_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _15294_/A VGND VGND VPWR VPWR _15387_/A sky130_fd_sc_hd__buf_2
XFILLER_8_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16722__B1 _16368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17033_ _17032_/Y VGND VGND VPWR VPWR _17074_/A sky130_fd_sc_hd__buf_2
XFILLER_172_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14245_ _14233_/A VGND VGND VPWR VPWR _14245_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_136_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23768_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_183_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14176_ _14176_/A VGND VGND VPWR VPWR _14176_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_199_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24666_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_152_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13127_ _24042_/Q _13127_/B VGND VGND VPWR VPWR _13145_/C sky130_fd_sc_hd__or2_4
XFILLER_97_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18984_ _18983_/Y _14674_/X _17430_/X _14674_/X VGND VGND VPWR VPWR _23907_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13058_ _13069_/A _13056_/X _13057_/X VGND VGND VPWR VPWR _25361_/D sky130_fd_sc_hd__and3_4
X_17935_ _17930_/A _17929_/Y _15922_/A VGND VGND VPWR VPWR _17935_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23220__B1 _22852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12009_ _12009_/A VGND VGND VPWR VPWR _12009_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13455__A _13423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15147__A2_N _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17866_ _17861_/A _17861_/B _17861_/D VGND VGND VPWR VPWR _17866_/X sky130_fd_sc_hd__or3_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16789__B1 _16537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16693__A1_N _16691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16817_ _16815_/Y _16816_/X _15732_/X _16816_/X VGND VGND VPWR VPWR _24445_/D sky130_fd_sc_hd__a2bb2o_4
X_19605_ _19605_/A VGND VGND VPWR VPWR _19605_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17797_ _17748_/X _17797_/B _17797_/C VGND VGND VPWR VPWR _17797_/X sky130_fd_sc_hd__and3_4
XANTENNA__13605__D _13786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19536_ _23713_/Q VGND VGND VPWR VPWR _21960_/B sky130_fd_sc_hd__inv_2
X_16748_ _16762_/A VGND VGND VPWR VPWR _16748_/X sky130_fd_sc_hd__buf_2
XFILLER_47_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17202__A1 _24636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17202__B2 _17263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19467_ _19465_/Y _19461_/X _19421_/X _19466_/X VGND VGND VPWR VPWR _23738_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _24504_/Q VGND VGND VPWR VPWR _16679_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24891__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ _18418_/A VGND VGND VPWR VPWR _18418_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19398_ _19396_/Y _19392_/X _19308_/X _19397_/X VGND VGND VPWR VPWR _23762_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24820__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18349_ _17461_/X _18349_/B VGND VGND VPWR VPWR _18352_/A sky130_fd_sc_hd__and2_4
XFILLER_159_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21360_ _21359_/X VGND VGND VPWR VPWR _21360_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_32_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_32_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20311_ _21933_/B _20308_/X _20000_/X _20308_/X VGND VGND VPWR VPWR _23440_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13527__B1 _13481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21291_ _21291_/A VGND VGND VPWR VPWR _21291_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22950__B _22946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23030_ _12825_/Y _21890_/X _16952_/Y _22839_/X VGND VGND VPWR VPWR _23030_/X sky130_fd_sc_hd__o22a_4
X_20242_ _23465_/Q VGND VGND VPWR VPWR _20242_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20273__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20173_ _20169_/Y _20172_/X _20102_/X _20172_/X VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18221__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_HCLK clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24981_ _24981_/CLK _15434_/Y HRESETn VGND VGND VPWR VPWR _15101_/A sky130_fd_sc_hd__dfrtp_4
X_23932_ _23475_/CLK _18918_/X VGND VGND VPWR VPWR _23932_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22678__A _22678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23863_ _23926_/CLK _23863_/D VGND VGND VPWR VPWR _23863_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22317__A2 _21312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22814_ _24601_/Q _23010_/B VGND VGND VPWR VPWR _22819_/B sky130_fd_sc_hd__or2_4
XFILLER_232_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23794_ _23794_/CLK _23794_/D VGND VGND VPWR VPWR _23794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_241_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24908__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25533_ _24386_/CLK _11839_/X HRESETn VGND VGND VPWR VPWR _25533_/Q sky130_fd_sc_hd__dfrtp_4
X_22745_ _22745_/A _22595_/B VGND VGND VPWR VPWR _22745_/X sky130_fd_sc_hd__and2_4
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22676_ _22294_/A _22676_/B _22676_/C _22675_/X VGND VGND VPWR VPWR _22676_/X sky130_fd_sc_hd__or4_4
X_25464_ _25456_/CLK _25464_/D HRESETn VGND VGND VPWR VPWR _12200_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24561__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21627_ _21646_/A _21625_/X _21626_/X VGND VGND VPWR VPWR _21627_/X sky130_fd_sc_hd__and3_4
X_24415_ _23577_/CLK _16882_/X HRESETn VGND VGND VPWR VPWR _24415_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23302__A _23302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25395_ _24812_/CLK _25395_/D HRESETn VGND VGND VPWR VPWR _25395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12360_ _12360_/A _12355_/X _12357_/X _12360_/D VGND VGND VPWR VPWR _12390_/A sky130_fd_sc_hd__or4_4
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21558_ _14496_/Y _21726_/B VGND VGND VPWR VPWR _21558_/X sky130_fd_sc_hd__or2_4
X_24346_ _24346_/CLK _24346_/D HRESETn VGND VGND VPWR VPWR _17251_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20509_ _20503_/X _20508_/Y VGND VGND VPWR VPWR _24092_/D sky130_fd_sc_hd__or2_4
XFILLER_166_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12291_ _12228_/Y _12212_/A _12288_/Y _12291_/D VGND VGND VPWR VPWR _12291_/X sky130_fd_sc_hd__or4_4
X_24277_ _24283_/CLK _24277_/D HRESETn VGND VGND VPWR VPWR _24277_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16180__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21489_ _18300_/B VGND VGND VPWR VPWR _21687_/A sky130_fd_sc_hd__buf_2
X_14030_ _14032_/B _14025_/Y _14026_/Y _14004_/A _14029_/Y VGND VGND VPWR VPWR _14030_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23228_ _23228_/A _22669_/B VGND VGND VPWR VPWR _23228_/X sky130_fd_sc_hd__or2_4
XFILLER_180_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_209_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24431_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_141_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20264__B1 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23159_ _22157_/C VGND VGND VPWR VPWR _23159_/X sky130_fd_sc_hd__buf_2
XFILLER_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15981_ _15974_/X _15977_/X _16248_/A _22644_/A _15975_/X VGND VGND VPWR VPWR _24765_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17720_ _24222_/Q _24221_/Q VGND VGND VPWR VPWR _17720_/X sky130_fd_sc_hd__and2_4
X_14932_ _25020_/Q _14931_/A _14930_/Y _14931_/Y VGND VGND VPWR VPWR _14933_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20139__A2_N _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22588__A _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ _17531_/Y _17651_/B VGND VGND VPWR VPWR _17652_/C sky130_fd_sc_hd__nand2_4
XFILLER_236_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14863_ _14854_/X _14862_/Y _24963_/Q _14854_/X VGND VGND VPWR VPWR _14863_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19709__B1 _19612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16586__A _24538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16602_ _16601_/Y _16597_/X _16248_/X _16597_/X VGND VGND VPWR VPWR _24532_/D sky130_fd_sc_hd__a2bb2o_4
X_13814_ _13811_/Y _13805_/X _13812_/X _13813_/X VGND VGND VPWR VPWR _25278_/D sky130_fd_sc_hd__a2bb2o_4
X_17582_ _17684_/A _17518_/Y _17522_/Y _17504_/Y VGND VGND VPWR VPWR _17589_/A sky130_fd_sc_hd__or4_4
XFILLER_35_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15994__A1 _15797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14794_ _14794_/A VGND VGND VPWR VPWR _17990_/A sky130_fd_sc_hd__inv_2
XFILLER_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22859__A3 _16468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19321_ _19320_/Y _19316_/X _19254_/X _19301_/Y VGND VGND VPWR VPWR _23789_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24649__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16533_ _16533_/A VGND VGND VPWR VPWR _16533_/X sky130_fd_sc_hd__buf_2
X_13745_ _13744_/X VGND VGND VPWR VPWR _19837_/A sky130_fd_sc_hd__buf_2
X_19252_ _19251_/Y _19249_/X _19184_/X _19249_/X VGND VGND VPWR VPWR _23814_/D sky130_fd_sc_hd__a2bb2o_4
X_16464_ _16464_/A _16464_/B _22754_/A _21173_/C VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__and4_4
XFILLER_189_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13676_ _13676_/A _20956_/A _20964_/A _20952_/A VGND VGND VPWR VPWR _13676_/X sky130_fd_sc_hd__or4_4
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20836__A _20836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18203_ _18107_/A _18203_/B _18203_/C VGND VGND VPWR VPWR _18203_/X sky130_fd_sc_hd__and3_4
X_15415_ _15415_/A _15399_/X VGND VGND VPWR VPWR _15417_/B sky130_fd_sc_hd__nand2_4
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23212__A _16662_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12627_ _12579_/Y _12574_/Y _12626_/X VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__or3_4
X_19183_ _19183_/A VGND VGND VPWR VPWR _19183_/Y sky130_fd_sc_hd__inv_2
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ HWDATA[27] VGND VGND VPWR VPWR _16395_/X sky130_fd_sc_hd__buf_2
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18134_ _18166_/A _18134_/B _18133_/X VGND VGND VPWR VPWR _18138_/B sky130_fd_sc_hd__and3_4
X_15346_ _15346_/A _15346_/B VGND VGND VPWR VPWR _15346_/X sky130_fd_sc_hd__or2_4
XFILLER_12_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12558_ _24869_/Q VGND VGND VPWR VPWR _12558_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13509__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18065_ _18199_/A _19195_/A VGND VGND VPWR VPWR _18067_/B sky130_fd_sc_hd__or2_4
X_15277_ _15259_/A _15280_/B _15183_/X VGND VGND VPWR VPWR _15277_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12354__A _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12489_ _12212_/X _12480_/X VGND VGND VPWR VPWR _12489_/X sky130_fd_sc_hd__or2_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17016_ _24398_/Q VGND VGND VPWR VPWR _17016_/Y sky130_fd_sc_hd__inv_2
X_14228_ _14228_/A VGND VGND VPWR VPWR _14229_/A sky130_fd_sc_hd__buf_2
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15665__A _15661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14159_ _14110_/A _14110_/B _14110_/A _14110_/B VGND VGND VPWR VPWR _14159_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18967_ _18965_/Y _18961_/X _17433_/X _18966_/X VGND VGND VPWR VPWR _23914_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17918_ _17905_/Y _17915_/A _17917_/X _22003_/A _17915_/Y VGND VGND VPWR VPWR _24260_/D
+ sky130_fd_sc_hd__a32o_4
X_18898_ _18876_/X _18890_/X _24124_/Q _24125_/Q _18893_/X VGND VGND VPWR VPWR _18898_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22498__A _21129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22952__C1 _22951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17849_ _17849_/A VGND VGND VPWR VPWR _17849_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20860_ _13667_/A _13667_/B _20859_/Y VGND VGND VPWR VPWR _20860_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19519_ _23719_/Q VGND VGND VPWR VPWR _21665_/B sky130_fd_sc_hd__inv_2
X_20791_ _20789_/Y _20785_/X _20790_/X VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22180__B1 _14137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22530_ _16706_/Y _22530_/B VGND VGND VPWR VPWR _22530_/X sky130_fd_sc_hd__and2_4
XANTENNA__18923__B2 _18922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16934__B1 _16164_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22461_ _15017_/Y _21085_/X _16468_/A _14925_/Y _22460_/X VGND VGND VPWR VPWR _22461_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_194_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21412_ _21412_/A _21410_/X _21411_/X VGND VGND VPWR VPWR _21412_/X sky130_fd_sc_hd__and3_4
X_24200_ _25145_/CLK _24200_/D HRESETn VGND VGND VPWR VPWR _18386_/A sky130_fd_sc_hd__dfrtp_4
X_25180_ _25181_/CLK _14325_/X HRESETn VGND VGND VPWR VPWR _25180_/Q sky130_fd_sc_hd__dfrtp_4
X_22392_ _22392_/A _20169_/Y VGND VGND VPWR VPWR _22392_/X sky130_fd_sc_hd__or2_4
XFILLER_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24131_ _24138_/CLK _24131_/D HRESETn VGND VGND VPWR VPWR _18686_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21343_ _21334_/Y VGND VGND VPWR VPWR _23148_/A sky130_fd_sc_hd__buf_2
XFILLER_163_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24062_ _24532_/CLK _20905_/X HRESETn VGND VGND VPWR VPWR _24062_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18439__B1 _16244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21274_ _21271_/A _20124_/Y VGND VGND VPWR VPWR _21275_/C sky130_fd_sc_hd__or2_4
XFILLER_162_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23013_ _23013_/A _23013_/B _23013_/C VGND VGND VPWR VPWR _23013_/X sky130_fd_sc_hd__and3_4
XANTENNA__20246__B1 _19753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20225_ _20225_/A VGND VGND VPWR VPWR _21622_/B sky130_fd_sc_hd__inv_2
XANTENNA__19047__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_182_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _23960_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_131_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20156_ _20150_/Y VGND VGND VPWR VPWR _20156_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_39_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _23597_/CLK sky130_fd_sc_hd__clkbuf_1
X_20087_ _20085_/Y _20081_/X _19772_/X _20086_/X VGND VGND VPWR VPWR _20087_/X sky130_fd_sc_hd__a2bb2o_4
X_24964_ _24339_/CLK _15469_/X HRESETn VGND VGND VPWR VPWR _13896_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23915_ _23913_/CLK _23915_/D VGND VGND VPWR VPWR _18963_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_217_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24895_ _24015_/CLK _15685_/X HRESETn VGND VGND VPWR VPWR _13680_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22201__A _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11860_ HWDATA[3] VGND VGND VPWR VPWR _11861_/A sky130_fd_sc_hd__buf_2
X_23846_ _24101_/CLK _19162_/X VGND VGND VPWR VPWR _19161_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24742__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _11789_/Y _11786_/X _11790_/X _11786_/X VGND VGND VPWR VPWR _25545_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_198_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20989_ _14131_/X _20988_/X _20996_/B VGND VGND VPWR VPWR _20989_/X sky130_fd_sc_hd__o21a_4
X_23777_ _23850_/CLK _19356_/X VGND VGND VPWR VPWR _18093_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12439__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22710__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _14299_/B VGND VGND VPWR VPWR _13533_/A sky130_fd_sc_hd__inv_2
X_25516_ _25520_/CLK _25516_/D HRESETn VGND VGND VPWR VPWR _25516_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22728_ _21714_/A _22724_/X _22728_/C VGND VGND VPWR VPWR _22728_/X sky130_fd_sc_hd__and3_4
XFILLER_198_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ _13257_/X _13461_/B VGND VGND VPWR VPWR _13461_/X sky130_fd_sc_hd__or2_4
X_25447_ _25443_/CLK _25447_/D HRESETn VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__dfrtp_4
X_22659_ _22643_/Y _22648_/Y _22656_/Y _21455_/X _22658_/X VGND VGND VPWR VPWR _22660_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_185_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15200_ _15199_/X VGND VGND VPWR VPWR _25039_/D sky130_fd_sc_hd__inv_2
X_12412_ _12401_/B _12401_/C _12411_/X _12408_/B VGND VGND VPWR VPWR _12412_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17030__A _17064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16180_ RsRx_S0 _16179_/Y _14781_/B VGND VGND VPWR VPWR _16180_/X sky130_fd_sc_hd__a21o_4
X_13392_ _13456_/A _13384_/X _13391_/X VGND VGND VPWR VPWR _13392_/X sky130_fd_sc_hd__and3_4
X_25378_ _25380_/CLK _25378_/D HRESETn VGND VGND VPWR VPWR _25378_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22871__A _22871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15131_ _24602_/Q VGND VGND VPWR VPWR _15131_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12343_ _24827_/Q VGND VGND VPWR VPWR _12343_/Y sky130_fd_sc_hd__inv_2
X_24329_ _23654_/CLK _24329_/D HRESETn VGND VGND VPWR VPWR _11657_/A sky130_fd_sc_hd__dfstp_4
XFILLER_166_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ _12273_/X _21715_/A _25439_/Q _12240_/Y VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__a2bb2o_4
X_15062_ _14910_/A _15060_/Y _25033_/Q _15061_/Y VGND VGND VPWR VPWR _15063_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21487__A _21679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20391__A _20385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14013_ _14013_/A _14013_/B _14010_/X _14022_/A VGND VGND VPWR VPWR _14014_/A sky130_fd_sc_hd__or4_4
X_19870_ _21917_/B _19867_/X _19800_/X _19867_/X VGND VGND VPWR VPWR _23601_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18821_ _18689_/B _18824_/B VGND VGND VPWR VPWR _18825_/B sky130_fd_sc_hd__or2_4
XFILLER_150_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18752_ _18752_/A _18751_/X VGND VGND VPWR VPWR _18753_/B sky130_fd_sc_hd__or2_4
XFILLER_191_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15964_ _12202_/Y _15962_/X _15963_/X _15962_/X VGND VGND VPWR VPWR _24774_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17703_ _17529_/Y _17703_/B VGND VGND VPWR VPWR _17704_/B sky130_fd_sc_hd__nand2_4
X_14915_ _14912_/X _14913_/Y _15195_/A _14914_/Y VGND VGND VPWR VPWR _14915_/X sky130_fd_sc_hd__a2bb2o_4
X_18683_ _18681_/Y _18683_/B VGND VGND VPWR VPWR _18701_/C sky130_fd_sc_hd__or2_4
XFILLER_248_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15895_ _15895_/A VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__buf_2
X_17634_ _17691_/A VGND VGND VPWR VPWR _17641_/A sky130_fd_sc_hd__buf_2
X_14846_ _14834_/X _14845_/Y _14826_/C _14834_/X VGND VGND VPWR VPWR _14846_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ _17691_/A VGND VGND VPWR VPWR _17598_/A sky130_fd_sc_hd__buf_2
XFILLER_63_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14777_ _14776_/X VGND VGND VPWR VPWR _14781_/B sky130_fd_sc_hd__inv_2
XANTENNA__15747__A1_N _12568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _11710_/A _11664_/A _11986_/X _11662_/A _11988_/X VGND VGND VPWR VPWR _11989_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17708__A2 _17610_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19304_ _23795_/Q VGND VGND VPWR VPWR _19304_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16515_/Y _16513_/X _16245_/X _16513_/X VGND VGND VPWR VPWR _16516_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13728_ _13697_/B _13716_/X _13727_/Y _13723_/X _11676_/A VGND VGND VPWR VPWR _13728_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_232_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17496_ _18335_/A _20079_/D _17494_/Y VGND VGND VPWR VPWR _17496_/X sky130_fd_sc_hd__a21o_4
X_19235_ _19234_/X VGND VGND VPWR VPWR _19249_/A sky130_fd_sc_hd__inv_2
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16447_ _16445_/Y _16442_/X _16364_/X _16446_/X VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__a2bb2o_4
X_13659_ _13659_/A _24067_/Q _13659_/C _13658_/X VGND VGND VPWR VPWR _20933_/B sky130_fd_sc_hd__or4_4
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23299__D _23298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19166_ _19166_/A _19166_/B _25079_/Q _13634_/X VGND VGND VPWR VPWR _19166_/X sky130_fd_sc_hd__or4_4
X_16378_ _16378_/A _16378_/B _16378_/C _16378_/D VGND VGND VPWR VPWR _16379_/A sky130_fd_sc_hd__or4_4
X_18117_ _18209_/A _18117_/B VGND VGND VPWR VPWR _18119_/B sky130_fd_sc_hd__or2_4
XFILLER_157_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15329_ _15302_/Y _15340_/A _15337_/A _15337_/B VGND VGND VPWR VPWR _15329_/X sky130_fd_sc_hd__or4_4
X_19097_ _23868_/Q VGND VGND VPWR VPWR _22379_/B sky130_fd_sc_hd__inv_2
XFILLER_144_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25144__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18048_ _18191_/A _18046_/X _18048_/C VGND VGND VPWR VPWR _18049_/C sky130_fd_sc_hd__and3_4
XFILLER_105_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19094__B1 _19048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20010_ _20010_/A VGND VGND VPWR VPWR _20010_/X sky130_fd_sc_hd__buf_2
XANTENNA__22005__B _20360_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_255_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _24979_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19999_ _23553_/Q VGND VGND VPWR VPWR _21956_/B sky130_fd_sc_hd__inv_2
XFILLER_247_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21961_ _21472_/A _21959_/X _21961_/C VGND VGND VPWR VPWR _21961_/X sky130_fd_sc_hd__and3_4
XFILLER_243_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23700_ _23716_/CLK _23700_/D VGND VGND VPWR VPWR _23700_/Q sky130_fd_sc_hd__dfxtp_4
X_20912_ _24064_/Q _20907_/X _20911_/X VGND VGND VPWR VPWR _20912_/Y sky130_fd_sc_hd__a21oi_4
X_21892_ _25442_/Q _23321_/A _21891_/X _21113_/X VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__a211o_4
X_24680_ _24657_/CLK _16206_/X HRESETn VGND VGND VPWR VPWR _23250_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _13660_/Y _13662_/B _13664_/B VGND VGND VPWR VPWR _20843_/X sky130_fd_sc_hd__o21a_4
X_23631_ _23631_/CLK _19781_/X VGND VGND VPWR VPWR _13403_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23350__C1 _23349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20774_ _20761_/X _20773_/Y _24915_/Q _20765_/X VGND VGND VPWR VPWR _24032_/D sky130_fd_sc_hd__a2bb2o_4
X_23562_ _23560_/CLK _19973_/X VGND VGND VPWR VPWR _19971_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25301_ _24233_/CLK _13706_/X HRESETn VGND VGND VPWR VPWR _25301_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22513_ _16524_/Y _22513_/B VGND VGND VPWR VPWR _22513_/X sky130_fd_sc_hd__and2_4
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23493_ _23493_/CLK _20168_/X VGND VGND VPWR VPWR _20167_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22444_ _21330_/X VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__buf_2
X_25232_ _25105_/CLK _25232_/D HRESETn VGND VGND VPWR VPWR _14042_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__14394__B1 _13844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22375_ _22394_/A _20211_/Y VGND VGND VPWR VPWR _22376_/C sky130_fd_sc_hd__or2_4
X_25163_ _24121_/CLK _14374_/X HRESETn VGND VGND VPWR VPWR _25163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21326_ _21293_/X _21304_/X _21308_/X _21319_/X _21325_/X VGND VGND VPWR VPWR _21326_/X
+ sky130_fd_sc_hd__o41a_4
X_24114_ _25145_/CLK _20979_/X HRESETn VGND VGND VPWR VPWR _12134_/B sky130_fd_sc_hd__dfrtp_4
X_25094_ _25093_/CLK _14609_/X HRESETn VGND VGND VPWR VPWR _25094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16905__A2_N _17767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21257_ _21257_/A _18933_/Y VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__or2_4
X_24045_ _24509_/CLK _20828_/X HRESETn VGND VGND VPWR VPWR _24045_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13818__A _13818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20208_ _21411_/B _20205_/X _20122_/X _20205_/X VGND VGND VPWR VPWR _23478_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18832__B1 _16510_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21188_ _21204_/A _21188_/B _21187_/X VGND VGND VPWR VPWR _21188_/X sky130_fd_sc_hd__and3_4
XFILLER_104_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15646__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20139_ _20138_/Y _20134_/X _20115_/X _20134_/X VGND VGND VPWR VPWR _23504_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ _12777_/X _12952_/X VGND VGND VPWR VPWR _12961_/X sky130_fd_sc_hd__or2_4
X_24947_ _23407_/CLK _15514_/X HRESETn VGND VGND VPWR VPWR _24947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14649__A _18051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19847__A2_N _19844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ _14687_/A VGND VGND VPWR VPWR _14700_/X sky130_fd_sc_hd__buf_2
X_11912_ _11883_/Y _11908_/Y _11895_/Y _11911_/X VGND VGND VPWR VPWR _11913_/A sky130_fd_sc_hd__a211o_4
XFILLER_85_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15680_ _21874_/A VGND VGND VPWR VPWR _22738_/A sky130_fd_sc_hd__buf_2
X_12892_ _12862_/X _12871_/X _12765_/Y VGND VGND VPWR VPWR _12893_/C sky130_fd_sc_hd__o21a_4
X_24878_ _24878_/CLK _15746_/X HRESETn VGND VGND VPWR VPWR _24878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_234_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16071__B1 _16070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ _14630_/X VGND VGND VPWR VPWR _14631_/Y sky130_fd_sc_hd__inv_2
X_11843_ _11840_/Y _11835_/X _11842_/X _11835_/X VGND VGND VPWR VPWR _11843_/X sky130_fd_sc_hd__a2bb2o_4
X_23829_ _23830_/CLK _23829_/D VGND VGND VPWR VPWR _18231_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17315_/X _17350_/B _17349_/X VGND VGND VPWR VPWR _17350_/X sky130_fd_sc_hd__and3_4
X_14562_ HREADY HSEL VGND VGND VPWR VPWR _14562_/Y sky130_fd_sc_hd__nand2_4
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11772_/Y _11769_/X _11773_/X _11769_/X VGND VGND VPWR VPWR _11774_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20386__A _20385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16300_/Y _16298_/X _15950_/X _16298_/X VGND VGND VPWR VPWR _24645_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13512_/Y _13510_/X _11847_/X _13510_/X VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _17270_/C _17278_/X _17271_/Y _17280_/X VGND VGND VPWR VPWR _17282_/A sky130_fd_sc_hd__a211o_4
XFILLER_201_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14493_ _21858_/A _14490_/X _14400_/X _14490_/X VGND VGND VPWR VPWR _14493_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14384__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19020_ _19020_/A VGND VGND VPWR VPWR _19020_/X sky130_fd_sc_hd__buf_2
X_16232_ _16231_/Y _16227_/X _15972_/X _16227_/X VGND VGND VPWR VPWR _24669_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13444_ _13153_/X _13444_/B _13444_/C VGND VGND VPWR VPWR _13448_/B sky130_fd_sc_hd__and3_4
XFILLER_173_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16163_ _16161_/Y _16162_/X _16070_/X _16162_/X VGND VGND VPWR VPWR _24692_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13375_ _13187_/X _13367_/X _13374_/X VGND VGND VPWR VPWR _13375_/X sky130_fd_sc_hd__and3_4
XFILLER_182_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15114_ _15114_/A VGND VGND VPWR VPWR _15114_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12326_ _25348_/Q VGND VGND VPWR VPWR _12326_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17874__A1 _17861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16094_ _22684_/B VGND VGND VPWR VPWR _22513_/B sky130_fd_sc_hd__buf_2
XFILLER_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12114__A1_N _12113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15045_ _14930_/Y VGND VGND VPWR VPWR _15259_/A sky130_fd_sc_hd__buf_2
X_19922_ _19921_/Y _19917_/X _19900_/X _19904_/Y VGND VGND VPWR VPWR _19922_/X sky130_fd_sc_hd__a2bb2o_4
X_12257_ _12257_/A VGND VGND VPWR VPWR _12294_/A sky130_fd_sc_hd__inv_2
XANTENNA__12699__B1 _12657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12188_ _12188_/A VGND VGND VPWR VPWR _12397_/A sky130_fd_sc_hd__inv_2
X_19853_ _19853_/A VGND VGND VPWR VPWR _19853_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15637__B1 _15636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20630__B1 _20680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18804_ _24140_/Q _18803_/Y VGND VGND VPWR VPWR _18806_/B sky130_fd_sc_hd__or2_4
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_22_0_HCLK clkbuf_8_23_0_HCLK/A VGND VGND VPWR VPWR _24327_/CLK sky130_fd_sc_hd__clkbuf_1
X_16996_ _16996_/A VGND VGND VPWR VPWR _16996_/Y sky130_fd_sc_hd__inv_2
X_19784_ _13467_/B VGND VGND VPWR VPWR _19784_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24664__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_85_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _25365_/CLK sky130_fd_sc_hd__clkbuf_1
X_15947_ _15947_/A VGND VGND VPWR VPWR _15947_/X sky130_fd_sc_hd__buf_2
X_18735_ _18683_/B _18735_/B VGND VGND VPWR VPWR _18736_/A sky130_fd_sc_hd__or2_4
XANTENNA__13463__A _13315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18666_ _16576_/A _18733_/A _16581_/Y _24151_/Q VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__a2bb2o_4
X_15878_ _12791_/Y _15877_/X _11758_/X _15877_/X VGND VGND VPWR VPWR _24819_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22776__A _22743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16062__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14829_ _14815_/C _14829_/B VGND VGND VPWR VPWR _14829_/Y sky130_fd_sc_hd__nor2_4
X_17617_ _17598_/A _17615_/X _17617_/C VGND VGND VPWR VPWR _24323_/D sky130_fd_sc_hd__and3_4
XFILLER_64_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18597_ _18425_/Y _18597_/B VGND VGND VPWR VPWR _18597_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22135__B1 _21565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17548_ _11782_/Y _17553_/A _25535_/Q _17585_/D VGND VGND VPWR VPWR _17548_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19000__B1 _18999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17479_ _20079_/D _18905_/D VGND VGND VPWR VPWR _17479_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19218_ _19216_/Y _19212_/X _19151_/X _19217_/X VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20490_ _14214_/A _20497_/B VGND VGND VPWR VPWR _20490_/X sky130_fd_sc_hd__or2_4
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19149_ _19147_/Y _19145_/X _19148_/X _19145_/X VGND VGND VPWR VPWR _23851_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22160_ _21043_/A _22159_/X _22144_/A _24830_/Q _15553_/X VGND VGND VPWR VPWR _22160_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_246_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21111_ _21058_/A _21104_/X _21111_/C VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__and3_4
XFILLER_160_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22091_ _22390_/A _22091_/B _22091_/C VGND VGND VPWR VPWR _22091_/X sky130_fd_sc_hd__and3_4
XFILLER_172_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21042_ _22533_/A VGND VGND VPWR VPWR _21042_/X sky130_fd_sc_hd__buf_2
XANTENNA__21855__A _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24801_ _24794_/CLK _15903_/X HRESETn VGND VGND VPWR VPWR _22605_/A sky130_fd_sc_hd__dfrtp_4
X_22993_ _21043_/A VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__buf_2
XANTENNA__24334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21716__A3 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24732_ _24732_/CLK _16057_/X HRESETn VGND VGND VPWR VPWR _24732_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_215_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21944_ _21948_/A _21944_/B VGND VGND VPWR VPWR _21945_/C sky130_fd_sc_hd__or2_4
XFILLER_216_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13804__C _13804_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _24169_/CLK _24663_/D HRESETn VGND VGND VPWR VPWR _24663_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ _16445_/A _23274_/B VGND VGND VPWR VPWR _21879_/B sky130_fd_sc_hd__or2_4
XFILLER_203_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23615_/CLK _19833_/X VGND VGND VPWR VPWR _23614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20822_/X VGND VGND VPWR VPWR _20826_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24594_ _24989_/CLK _16439_/X HRESETn VGND VGND VPWR VPWR _15121_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_202_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23684_/CLK _23545_/D VGND VGND VPWR VPWR _20024_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20757_ _20753_/X VGND VGND VPWR VPWR _20757_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22429__A1 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20688_ _20683_/X _20687_/X _20621_/B VGND VGND VPWR VPWR _20688_/X sky130_fd_sc_hd__o21a_4
X_23476_ _23475_/CLK _20215_/X VGND VGND VPWR VPWR _20211_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_195_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25215_ _25215_/CLK _14193_/Y HRESETn VGND VGND VPWR VPWR _14190_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_183_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22427_ _21604_/A _22427_/B VGND VGND VPWR VPWR _22427_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13160_ _13271_/A VGND VGND VPWR VPWR _13443_/A sky130_fd_sc_hd__buf_2
X_25146_ _25223_/CLK _14433_/X HRESETn VGND VGND VPWR VPWR _25146_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22358_ _22032_/A _22358_/B VGND VGND VPWR VPWR _22358_/X sky130_fd_sc_hd__or2_4
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12111_ _12123_/A VGND VGND VPWR VPWR _12111_/X sky130_fd_sc_hd__buf_2
X_13091_ _12351_/Y _13091_/B VGND VGND VPWR VPWR _13107_/B sky130_fd_sc_hd__or2_4
X_21309_ _21872_/A VGND VGND VPWR VPWR _22723_/A sky130_fd_sc_hd__buf_2
X_22289_ _22289_/A VGND VGND VPWR VPWR _22289_/X sky130_fd_sc_hd__buf_2
X_25077_ _25077_/CLK _25077_/D HRESETn VGND VGND VPWR VPWR _13626_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12042_ _25498_/Q VGND VGND VPWR VPWR _12042_/Y sky130_fd_sc_hd__inv_2
X_24028_ _24495_/CLK _20755_/X HRESETn VGND VGND VPWR VPWR _20752_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15882__A3 _15732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15619__B1 _11827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16850_ _14943_/Y _16846_/X _16609_/X _16849_/X VGND VGND VPWR VPWR _16850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15801_ _15826_/A VGND VGND VPWR VPWR _15802_/A sky130_fd_sc_hd__buf_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16292__B1 _11752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16781_ _15032_/Y _16779_/X _11830_/X _16779_/X VGND VGND VPWR VPWR _24461_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13993_ _14053_/C _14028_/D _14027_/C _14027_/D VGND VGND VPWR VPWR _13993_/X sky130_fd_sc_hd__and4_4
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18520_ _18517_/A _18517_/B VGND VGND VPWR VPWR _18521_/C sky130_fd_sc_hd__nand2_4
XFILLER_234_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13283__A _13322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22904__A2 _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15732_ HWDATA[26] VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__buf_2
X_12944_ _22678_/A _12944_/B VGND VGND VPWR VPWR _12945_/C sky130_fd_sc_hd__or2_4
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18451_ _18451_/A _18451_/B _18451_/C _18451_/D VGND VGND VPWR VPWR _18451_/X sky130_fd_sc_hd__or4_4
X_15663_ _15662_/Y VGND VGND VPWR VPWR _15663_/X sky130_fd_sc_hd__buf_2
XFILLER_206_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12875_ _12908_/A VGND VGND VPWR VPWR _12875_/X sky130_fd_sc_hd__buf_2
XFILLER_233_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17402_ _17402_/A _17402_/B VGND VGND VPWR VPWR _20653_/A sky130_fd_sc_hd__or2_4
XPHY_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14610_/B _14613_/Y _14608_/X _14611_/X _25092_/Q VGND VGND VPWR VPWR _14614_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ HWDATA[11] VGND VGND VPWR VPWR _16252_/A sky130_fd_sc_hd__buf_2
X_18382_ _18381_/Y _18379_/X _24201_/Q _18379_/X VGND VGND VPWR VPWR _24202_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15594_/A VGND VGND VPWR VPWR _23003_/A sky130_fd_sc_hd__inv_2
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17330_/B VGND VGND VPWR VPWR _17333_/Y sky130_fd_sc_hd__inv_2
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14545_/A VGND VGND VPWR VPWR _14545_/Y sky130_fd_sc_hd__inv_2
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _25554_/Q VGND VGND VPWR VPWR _11757_/Y sky130_fd_sc_hd__inv_2
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17264_ _17257_/Y _17258_/Y _17261_/X _17318_/A VGND VGND VPWR VPWR _17265_/B sky130_fd_sc_hd__or4_4
X_14476_ _14474_/Y _14475_/X _14404_/X _14475_/X VGND VGND VPWR VPWR _14476_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _11688_/A VGND VGND VPWR VPWR _11688_/Y sky130_fd_sc_hd__inv_2
X_19003_ _19002_/X VGND VGND VPWR VPWR _19020_/A sky130_fd_sc_hd__inv_2
X_16215_ _16227_/A VGND VGND VPWR VPWR _16215_/X sky130_fd_sc_hd__buf_2
X_13427_ _13322_/A _13425_/X _13426_/X VGND VGND VPWR VPWR _13427_/X sky130_fd_sc_hd__and3_4
XANTENNA__15938__A _15796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17195_ _17195_/A VGND VGND VPWR VPWR _17248_/B sky130_fd_sc_hd__inv_2
XFILLER_155_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16146_ _16145_/Y _16141_/X _11822_/X _16141_/X VGND VGND VPWR VPWR _16146_/X sky130_fd_sc_hd__a2bb2o_4
X_13358_ _13454_/A _13358_/B _13357_/X VGND VGND VPWR VPWR _13359_/C sky130_fd_sc_hd__and3_4
XANTENNA__22840__A1 _12819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12309_ _12308_/Y _24850_/Q _12308_/Y _24850_/Q VGND VGND VPWR VPWR _12310_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13458__A _13282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19049__B1 _19048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16077_ _16075_/Y _16069_/X _15480_/X _16076_/X VGND VGND VPWR VPWR _16077_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13289_ _13242_/X _13287_/X _13289_/C VGND VGND VPWR VPWR _13289_/X sky130_fd_sc_hd__and3_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24845__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15028_ _24464_/Q VGND VGND VPWR VPWR _22682_/A sky130_fd_sc_hd__inv_2
X_19905_ _19904_/Y VGND VGND VPWR VPWR _19905_/X sky130_fd_sc_hd__buf_2
XANTENNA__21675__A _21675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15873__A3 _15562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19836_ _23612_/Q VGND VGND VPWR VPWR _22371_/B sky130_fd_sc_hd__inv_2
XANTENNA__19145__A _19159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16283__B1 _24650_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _19763_/Y _19766_/X _19677_/X _19766_/X VGND VGND VPWR VPWR _19767_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13097__B1 _13040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16979_ _16084_/Y _24378_/Q _16084_/Y _24378_/Q VGND VGND VPWR VPWR _16979_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21159__B2 _14442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22184__A1_N _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18718_ _18720_/B VGND VGND VPWR VPWR _18719_/B sky130_fd_sc_hd__inv_2
XANTENNA__19221__B1 _19220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19698_ _19698_/A VGND VGND VPWR VPWR _19698_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18649_ _24521_/Q _18689_/C _16620_/A _18809_/A VGND VGND VPWR VPWR _18649_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_240_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17783__B1 _16964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21660_ _13789_/X VGND VGND VPWR VPWR _21660_/X sky130_fd_sc_hd__buf_2
XANTENNA__22659__B2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20611_ _20448_/X _20609_/X _20610_/Y VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__and3_4
X_21591_ _21591_/A VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__buf_2
X_20542_ _20540_/B _20537_/B _20508_/Y _20541_/X VGND VGND VPWR VPWR _24084_/D sky130_fd_sc_hd__a211o_4
X_23330_ _22677_/B _23327_/Y _23168_/X _23329_/X VGND VGND VPWR VPWR _23330_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20473_ _14082_/A _20473_/B VGND VGND VPWR VPWR _20476_/C sky130_fd_sc_hd__and2_4
X_23261_ _16474_/A _23087_/B _22954_/C VGND VGND VPWR VPWR _23261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15848__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25000_ _24989_/CLK _15373_/X HRESETn VGND VGND VPWR VPWR _25000_/Q sky130_fd_sc_hd__dfrtp_4
X_22212_ _22227_/A _20104_/Y VGND VGND VPWR VPWR _22212_/X sky130_fd_sc_hd__or2_4
X_23192_ _24445_/Q _22947_/X _23015_/X _23191_/X VGND VGND VPWR VPWR _23192_/X sky130_fd_sc_hd__a211o_4
XFILLER_180_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22831__A1 _24537_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15849__B1 _15848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22143_ _21300_/Y VGND VGND VPWR VPWR _22144_/A sky130_fd_sc_hd__buf_2
XFILLER_161_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25200__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24586__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22074_ _22095_/A _20218_/Y VGND VGND VPWR VPWR _22075_/C sky130_fd_sc_hd__or2_4
XFILLER_161_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _21130_/A _21025_/B VGND VGND VPWR VPWR _21025_/X sky130_fd_sc_hd__and2_4
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16274__B1 _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20070__B2 _20065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24111__D MSI_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14199__A _14199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12835__B1 _12834_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22976_ _22771_/X _22974_/X _22702_/X _22975_/X VGND VGND VPWR VPWR _22976_/X sky130_fd_sc_hd__o22a_4
XFILLER_228_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24715_ _24715_/CLK _24715_/D HRESETn VGND VGND VPWR VPWR _24715_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21927_ _21923_/X _21926_/X _22221_/A VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__o21a_4
XFILLER_215_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12660_ _12660_/A _12660_/B VGND VGND VPWR VPWR _12669_/B sky130_fd_sc_hd__or2_4
X_24646_ _24639_/CLK _24646_/D HRESETn VGND VGND VPWR VPWR _16296_/A sky130_fd_sc_hd__dfrtp_4
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _21858_/A _21726_/B VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__or2_4
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23311__A2 _22485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20809_/A VGND VGND VPWR VPWR _20809_/Y sky130_fd_sc_hd__inv_2
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12591_/A VGND VGND VPWR VPWR _12591_/Y sky130_fd_sc_hd__inv_2
X_24577_ _24562_/CLK _16486_/X HRESETn VGND VGND VPWR VPWR _24577_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17526__B1 _11757_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21789_ _22387_/A _21787_/X _21788_/X VGND VGND VPWR VPWR _21789_/X sky130_fd_sc_hd__and3_4
XANTENNA__25303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _25177_/Q _14308_/Y _25176_/Q _14316_/A VGND VGND VPWR VPWR _14330_/X sky130_fd_sc_hd__o22a_4
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23528_ _23513_/CLK _23528_/D VGND VGND VPWR VPWR _23528_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _24009_/Q _14257_/X _14260_/X VGND VGND VPWR VPWR _14261_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23459_ _23459_/CLK _23459_/D VGND VGND VPWR VPWR _20260_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19080__A2_N _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ _14385_/A _16378_/B _16378_/C _15791_/D VGND VGND VPWR VPWR _16000_/X sky130_fd_sc_hd__or4_4
X_13212_ _13212_/A VGND VGND VPWR VPWR _13417_/A sky130_fd_sc_hd__buf_2
X_14192_ _14181_/X _14190_/Y _14138_/X _14191_/Y _14141_/A VGND VGND VPWR VPWR _14192_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ _20797_/A _20794_/B _13143_/C VGND VGND VPWR VPWR _13143_/X sky130_fd_sc_hd__or3_4
X_25129_ _25154_/CLK _14476_/X HRESETn VGND VGND VPWR VPWR _14474_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17973__A _17973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23357__A2_N _21834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21495__A _21687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13074_ _13074_/A VGND VGND VPWR VPWR _13074_/Y sky130_fd_sc_hd__inv_2
X_17951_ _17951_/A _17951_/B VGND VGND VPWR VPWR _17952_/C sky130_fd_sc_hd__or2_4
XANTENNA__15855__A3 _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12025_ _12024_/X VGND VGND VPWR VPWR _12025_/Y sky130_fd_sc_hd__inv_2
X_16902_ _22201_/A _16901_/Y _16108_/Y _16910_/A VGND VGND VPWR VPWR _16904_/C sky130_fd_sc_hd__a2bb2o_4
X_17882_ _17860_/D VGND VGND VPWR VPWR _17883_/B sky130_fd_sc_hd__inv_2
XFILLER_39_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_30_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16265__B1 _16070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19621_ _19619_/Y _19615_/X _19620_/X _19615_/A VGND VGND VPWR VPWR _19621_/X sky130_fd_sc_hd__a2bb2o_4
X_16833_ _16857_/A VGND VGND VPWR VPWR _16853_/A sky130_fd_sc_hd__buf_2
X_16764_ _16764_/A VGND VGND VPWR VPWR _16764_/Y sky130_fd_sc_hd__inv_2
X_19552_ _19565_/A VGND VGND VPWR VPWR _19552_/X sky130_fd_sc_hd__buf_2
X_13976_ _13976_/A VGND VGND VPWR VPWR _13976_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16017__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15715_ _21172_/B VGND VGND VPWR VPWR _15715_/X sky130_fd_sc_hd__buf_2
X_18503_ _18488_/A _18710_/A VGND VGND VPWR VPWR _18503_/X sky130_fd_sc_hd__and2_4
X_12927_ _12927_/A _12927_/B _12926_/Y VGND VGND VPWR VPWR _25391_/D sky130_fd_sc_hd__and3_4
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16695_ _16694_/Y _16692_/X _15754_/X _16692_/X VGND VGND VPWR VPWR _16695_/X sky130_fd_sc_hd__a2bb2o_4
X_19483_ _19483_/A VGND VGND VPWR VPWR _19483_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_159_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _25145_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_206_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15646_ _15645_/Y _15641_/X _14479_/X _15641_/X VGND VGND VPWR VPWR _24899_/D sky130_fd_sc_hd__a2bb2o_4
X_18434_ _18434_/A VGND VGND VPWR VPWR _18482_/A sky130_fd_sc_hd__inv_2
X_12858_ _12822_/A _12858_/B _12857_/Y _12834_/Y VGND VGND VPWR VPWR _12858_/X sky130_fd_sc_hd__or4_4
XFILLER_179_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _16238_/A VGND VGND VPWR VPWR _11809_/X sky130_fd_sc_hd__buf_2
X_18365_ _18364_/X VGND VGND VPWR VPWR _18365_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12054__A1 _24111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15577_ _15584_/A VGND VGND VPWR VPWR _15577_/X sky130_fd_sc_hd__buf_2
XFILLER_159_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12789_ _25392_/Q _22913_/A _12787_/Y _12788_/Y VGND VGND VPWR VPWR _12799_/A sky130_fd_sc_hd__o22a_4
XANTENNA__25044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17257_/Y _17258_/Y _17355_/B _17256_/X VGND VGND VPWR VPWR _17317_/C sky130_fd_sc_hd__or4_4
XFILLER_175_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14528_ _25113_/Q _14520_/X _25112_/Q _14522_/X VGND VGND VPWR VPWR _14528_/X sky130_fd_sc_hd__o22a_4
X_18296_ _17723_/X _17713_/X _18294_/X VGND VGND VPWR VPWR _18296_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21864__A2 _12107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17247_ _24371_/Q VGND VGND VPWR VPWR _17305_/A sky130_fd_sc_hd__inv_2
X_14459_ _14186_/Y _14457_/X _14248_/X _14457_/X VGND VGND VPWR VPWR _25136_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23066__B2 _22924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17178_ _17178_/A VGND VGND VPWR VPWR _17378_/A sky130_fd_sc_hd__buf_2
XFILLER_115_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16129_ _16127_/Y _16123_/X _15967_/X _16128_/X VGND VGND VPWR VPWR _24705_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15846__A3 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19442__B1 _19418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19819_ _19819_/A VGND VGND VPWR VPWR _19819_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22830_ _24569_/Q _22954_/B _22830_/C VGND VGND VPWR VPWR _22830_/X sky130_fd_sc_hd__and3_4
XANTENNA__23979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_55_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22761_ _21307_/B _22760_/X _21314_/X _24736_/Q _21317_/X VGND VGND VPWR VPWR _22761_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_25_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21552__A1 _21547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18219__A _18059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21552__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24500_ _24500_/CLK _16690_/X HRESETn VGND VGND VPWR VPWR _16689_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_213_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21712_ _21712_/A _23016_/A VGND VGND VPWR VPWR _21712_/X sky130_fd_sc_hd__or2_4
X_25480_ _24196_/CLK _25480_/D HRESETn VGND VGND VPWR VPWR _25480_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16246__A1_N _16244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22692_ _21113_/X _22690_/X _22468_/X _22691_/X VGND VGND VPWR VPWR _22692_/X sky130_fd_sc_hd__o22a_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21290__D _21290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _24431_/CLK _24431_/D HRESETn VGND VGND VPWR VPWR _16843_/A sky130_fd_sc_hd__dfrtp_4
X_21643_ _21637_/X _21642_/X _14721_/X VGND VGND VPWR VPWR _21651_/B sky130_fd_sc_hd__o21a_4
XFILLER_178_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24362_ _24346_/CLK _24362_/D HRESETn VGND VGND VPWR VPWR _17262_/A sky130_fd_sc_hd__dfrtp_4
X_21574_ _21574_/A VGND VGND VPWR VPWR _21741_/A sky130_fd_sc_hd__buf_2
X_23313_ _16387_/A _23313_/B VGND VGND VPWR VPWR _23313_/X sky130_fd_sc_hd__or2_4
X_20525_ _20525_/A _20525_/B _20504_/A _20511_/C VGND VGND VPWR VPWR _20525_/X sky130_fd_sc_hd__and4_4
X_24293_ _24272_/CLK _17784_/Y HRESETn VGND VGND VPWR VPWR _24293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24767__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20456_ _14073_/A _20443_/X _20447_/Y _20455_/X VGND VGND VPWR VPWR _20456_/X sky130_fd_sc_hd__a211o_4
X_23244_ _23244_/A _23303_/B VGND VGND VPWR VPWR _23244_/X sky130_fd_sc_hd__and2_4
X_20387_ _22364_/B _20386_/X _19626_/A _20386_/X VGND VGND VPWR VPWR _23411_/D sky130_fd_sc_hd__a2bb2o_4
X_23175_ _17245_/Y _22926_/X _25399_/Q _22927_/X VGND VGND VPWR VPWR _23176_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22126_ _12120_/Y _21579_/X _18383_/Y _21580_/X VGND VGND VPWR VPWR _22126_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22057_ _14734_/A _19614_/Y _22054_/X _22056_/X VGND VGND VPWR VPWR _22058_/A sky130_fd_sc_hd__o22a_4
XFILLER_247_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12730__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23019__B _23014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21008_ _21008_/A _21008_/B VGND VGND VPWR VPWR _21008_/X sky130_fd_sc_hd__and2_4
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13830_ _13848_/A VGND VGND VPWR VPWR _13838_/A sky130_fd_sc_hd__buf_2
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21762__B _21746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25555__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13761_ _13760_/X VGND VGND VPWR VPWR _13761_/X sky130_fd_sc_hd__buf_2
XFILLER_244_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11784__A1_N _11782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22959_ _24741_/Q _21039_/X _21068_/X _22958_/X VGND VGND VPWR VPWR _22960_/C sky130_fd_sc_hd__a211o_4
XFILLER_16_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15500_ _15503_/A VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__buf_2
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12712_ _12590_/Y _12712_/B VGND VGND VPWR VPWR _12732_/A sky130_fd_sc_hd__or2_4
X_16480_ _24579_/Q VGND VGND VPWR VPWR _16480_/Y sky130_fd_sc_hd__inv_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _13736_/A _13691_/X VGND VGND VPWR VPWR _13692_/X sky130_fd_sc_hd__or2_4
XFILLER_204_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15431_ _15311_/A _15430_/Y VGND VGND VPWR VPWR _15432_/B sky130_fd_sc_hd__or2_4
X_12643_ _12642_/X VGND VGND VPWR VPWR _12644_/B sky130_fd_sc_hd__inv_2
X_24629_ _24629_/CLK _24629_/D HRESETn VGND VGND VPWR VPWR _24629_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18150_ _17979_/A _18150_/B VGND VGND VPWR VPWR _18150_/X sky130_fd_sc_hd__or2_4
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15362_ _15362_/A _15361_/X VGND VGND VPWR VPWR _15363_/A sky130_fd_sc_hd__or2_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _12574_/A VGND VGND VPWR VPWR _12574_/Y sky130_fd_sc_hd__inv_2
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21846__A2 _21844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _17044_/C _17101_/B VGND VGND VPWR VPWR _17101_/X sky130_fd_sc_hd__or2_4
XANTENNA__11795__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _14313_/A VGND VGND VPWR VPWR _14313_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18081_ _18178_/A _18081_/B VGND VGND VPWR VPWR _18082_/C sky130_fd_sc_hd__or2_4
XFILLER_8_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _15293_/A _15293_/B _15292_/Y VGND VGND VPWR VPWR _25014_/D sky130_fd_sc_hd__and3_4
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12905__A _12817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17032_ _24650_/Q VGND VGND VPWR VPWR _17032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21059__B1 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14244_ _25201_/Q VGND VGND VPWR VPWR _14244_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14733__B1 _13748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14175_ _14131_/X _14108_/B _14107_/D _14174_/X VGND VGND VPWR VPWR _14176_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19672__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16486__B1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13126_ _13126_/A VGND VGND VPWR VPWR _13126_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18983_ _23907_/Q VGND VGND VPWR VPWR _18983_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _12996_/Y _13055_/A VGND VGND VPWR VPWR _13057_/X sky130_fd_sc_hd__or2_4
X_17934_ _17933_/X VGND VGND VPWR VPWR _17934_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12008_ _20971_/A _12000_/B _12007_/Y VGND VGND VPWR VPWR _12010_/A sky130_fd_sc_hd__o21a_4
XFILLER_239_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17865_ _17881_/A _17865_/B _17865_/C VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__and3_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19604_ _19603_/Y _19601_/X _19418_/X _19601_/X VGND VGND VPWR VPWR _23691_/D sky130_fd_sc_hd__a2bb2o_4
X_16816_ _16810_/X VGND VGND VPWR VPWR _16816_/X sky130_fd_sc_hd__buf_2
XFILLER_94_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12374__A2_N _24829_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17796_ _16910_/Y _17793_/X VGND VGND VPWR VPWR _17797_/C sky130_fd_sc_hd__or2_4
XFILLER_93_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19535_ _22039_/B _19529_/X _11948_/X _19534_/X VGND VGND VPWR VPWR _19535_/X sky130_fd_sc_hd__a2bb2o_4
X_13959_ _13949_/Y _13953_/Y _13956_/Y _13958_/X VGND VGND VPWR VPWR _13959_/X sky130_fd_sc_hd__or4_4
X_16747_ _15024_/Y _16743_/X _16395_/X _16743_/X VGND VGND VPWR VPWR _24478_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22731__B1 _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13471__A _13186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16678_ _16677_/Y _16673_/X _16410_/X _16673_/X VGND VGND VPWR VPWR _24505_/D sky130_fd_sc_hd__a2bb2o_4
X_19466_ _19460_/Y VGND VGND VPWR VPWR _19466_/X sky130_fd_sc_hd__buf_2
XFILLER_179_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22784__A _21436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18417_ _16214_/A _24187_/Q _16214_/Y _18517_/A VGND VGND VPWR VPWR _18420_/C sky130_fd_sc_hd__o22a_4
X_15629_ _14420_/A VGND VGND VPWR VPWR _15629_/X sky130_fd_sc_hd__buf_2
XFILLER_50_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19397_ _19391_/X VGND VGND VPWR VPWR _19397_/X sky130_fd_sc_hd__buf_2
XFILLER_210_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18348_ _13285_/A _18347_/X _13285_/A _18347_/X VGND VGND VPWR VPWR _18348_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18279_ _18278_/X _20405_/A VGND VGND VPWR VPWR _18279_/X sky130_fd_sc_hd__or2_4
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20310_ _23440_/Q VGND VGND VPWR VPWR _21933_/B sky130_fd_sc_hd__inv_2
XANTENNA__24860__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21290_ _21290_/A _21226_/X _21290_/C _21290_/D VGND VGND VPWR VPWR _21291_/A sky130_fd_sc_hd__and4_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12735__C1 _12662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22798__B1 _25389_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20241_ _20239_/Y _20235_/X _19772_/X _20240_/X VGND VGND VPWR VPWR _23466_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19663__B1 _19560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16477__B1 _16389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20172_ _20172_/A VGND VGND VPWR VPWR _20172_/X sky130_fd_sc_hd__buf_2
XANTENNA__12750__A2 _12403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24980_ _24979_/CLK _15445_/Y HRESETn VGND VGND VPWR VPWR _24980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16170__A1_N _16169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23931_ _23475_/CLK _18920_/X VGND VGND VPWR VPWR _23931_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22678__B _22678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23862_ _25066_/CLK _23862_/D VGND VGND VPWR VPWR _23862_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22813_ _22813_/A VGND VGND VPWR VPWR _23020_/A sky130_fd_sc_hd__buf_2
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23793_ _23794_/CLK _19312_/X VGND VGND VPWR VPWR _23793_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_226_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22722__B1 _21121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25532_ _24386_/CLK _11843_/X HRESETn VGND VGND VPWR VPWR _25532_/Q sky130_fd_sc_hd__dfrtp_4
X_22744_ _13564_/Y _22706_/B VGND VGND VPWR VPWR _22744_/X sky130_fd_sc_hd__and2_4
XFILLER_241_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16401__B1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_142_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _23794_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_197_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25463_ _25380_/CLK _12429_/X HRESETn VGND VGND VPWR VPWR _25463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17788__A _16925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22675_ _22678_/B _22671_/Y _21079_/A _22674_/X VGND VGND VPWR VPWR _22675_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24414_ _23529_/CLK _24414_/D HRESETn VGND VGND VPWR VPWR _20115_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21289__B1 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21626_ _21629_/A _21626_/B VGND VGND VPWR VPWR _21626_/X sky130_fd_sc_hd__or2_4
X_25394_ _25392_/CLK _25394_/D HRESETn VGND VGND VPWR VPWR _12857_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24345_ _24343_/CLK _24345_/D HRESETn VGND VGND VPWR VPWR _21010_/A sky130_fd_sc_hd__dfstp_4
X_21557_ _21293_/X _21534_/X _21540_/X _21553_/X _21556_/X VGND VGND VPWR VPWR _21557_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20508_ _13982_/A _20508_/B VGND VGND VPWR VPWR _20508_/Y sky130_fd_sc_hd__nor2_4
X_12290_ _12290_/A _12232_/Y _12513_/A VGND VGND VPWR VPWR _12291_/D sky130_fd_sc_hd__or3_4
X_24276_ _24283_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _17762_/A sky130_fd_sc_hd__dfrtp_4
X_21488_ _17716_/A VGND VGND VPWR VPWR _21493_/A sky130_fd_sc_hd__buf_2
XFILLER_180_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23227_ _23208_/X _23211_/X _23215_/Y _23226_/X VGND VGND VPWR VPWR HRDATA[27] sky130_fd_sc_hd__a211o_4
X_20439_ _20438_/X VGND VGND VPWR VPWR _23938_/D sky130_fd_sc_hd__buf_2
XANTENNA__19654__B1 _19439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23158_ _24779_/Q _23158_/B VGND VGND VPWR VPWR _23158_/X sky130_fd_sc_hd__or2_4
XFILLER_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22109_ _24557_/Q _21069_/B _21344_/X VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__o21a_4
XFILLER_164_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17028__A _17355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15980_ _15974_/X _15977_/X _16245_/A _22665_/A _15975_/X VGND VGND VPWR VPWR _24766_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23089_ _23025_/A _23089_/B _23088_/X VGND VGND VPWR VPWR _23089_/X sky130_fd_sc_hd__and3_4
X_14931_ _14931_/A VGND VGND VPWR VPWR _14931_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21773__A _14761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22961__B1 _16950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14862_ _14862_/A VGND VGND VPWR VPWR _14862_/Y sky130_fd_sc_hd__inv_2
X_17650_ _17578_/B _17649_/X VGND VGND VPWR VPWR _17651_/B sky130_fd_sc_hd__or2_4
XFILLER_235_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13813_ _13805_/A VGND VGND VPWR VPWR _13813_/X sky130_fd_sc_hd__buf_2
X_16601_ _16601_/A VGND VGND VPWR VPWR _16601_/Y sky130_fd_sc_hd__inv_2
X_17581_ _17581_/A VGND VGND VPWR VPWR _17581_/Y sky130_fd_sc_hd__inv_2
X_14793_ _14785_/A _14791_/X _14792_/Y VGND VGND VPWR VPWR _14793_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15994__A2 _15895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16532_ _16532_/A VGND VGND VPWR VPWR _16532_/Y sky130_fd_sc_hd__inv_2
X_19320_ _13460_/B VGND VGND VPWR VPWR _19320_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13744_ _13744_/A VGND VGND VPWR VPWR _13744_/X sky130_fd_sc_hd__buf_2
XFILLER_188_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16463_ _16462_/X VGND VGND VPWR VPWR _21173_/C sky130_fd_sc_hd__inv_2
X_19251_ _13413_/B VGND VGND VPWR VPWR _19251_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13675_ _20944_/A _20944_/B _13675_/C _13674_/X VGND VGND VPWR VPWR _20952_/A sky130_fd_sc_hd__or4_4
XFILLER_204_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16943__B2 _17751_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15414_ _15393_/A _15401_/X _15413_/Y VGND VGND VPWR VPWR _24988_/D sky130_fd_sc_hd__and3_4
X_18202_ _18138_/A _18202_/B _18202_/C VGND VGND VPWR VPWR _18203_/C sky130_fd_sc_hd__or3_4
XANTENNA__24689__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12626_ _12621_/X _12623_/X _12626_/C VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__or3_4
X_19182_ _19180_/Y _19181_/X _19091_/X _19181_/X VGND VGND VPWR VPWR _19182_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ _15154_/Y _16391_/X _16393_/X _16391_/X VGND VGND VPWR VPWR _24613_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23212__B _23303_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ _18165_/A _18133_/B VGND VGND VPWR VPWR _18133_/X sky130_fd_sc_hd__or2_4
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24618__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15345_ _15388_/A _15314_/X _15345_/C _15307_/X VGND VGND VPWR VPWR _15346_/B sky130_fd_sc_hd__or4_4
X_12557_ _12557_/A VGND VGND VPWR VPWR _12621_/A sky130_fd_sc_hd__inv_2
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15011__A _15011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18064_ _18098_/A VGND VGND VPWR VPWR _18199_/A sky130_fd_sc_hd__buf_2
X_15276_ _15276_/A _15276_/B VGND VGND VPWR VPWR _15280_/B sky130_fd_sc_hd__or2_4
X_12488_ _12488_/A VGND VGND VPWR VPWR _12488_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20231__A2_N _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17015_ _16075_/Y _17051_/A _24749_/Q _17034_/A VGND VGND VPWR VPWR _17015_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14227_ _14227_/A VGND VGND VPWR VPWR _14227_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19418__A _19148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14158_ _14155_/X _14157_/Y _25144_/Q _14155_/X VGND VGND VPWR VPWR _14158_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13109_ _13092_/X _13107_/Y _13121_/C VGND VGND VPWR VPWR _13109_/X sky130_fd_sc_hd__and3_4
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13466__A _13217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14089_ _24011_/Q _14078_/X _14082_/X _13999_/C _14085_/X VGND VGND VPWR VPWR _14089_/X
+ sky130_fd_sc_hd__a32o_4
X_18966_ _18974_/A VGND VGND VPWR VPWR _18966_/X sky130_fd_sc_hd__buf_2
XFILLER_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22779__A _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17917_ _22005_/A _17904_/X VGND VGND VPWR VPWR _17917_/X sky130_fd_sc_hd__or2_4
X_18897_ _18876_/X _18890_/X _24125_/Q _24126_/Q _18893_/X VGND VGND VPWR VPWR _24126_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17848_ _17763_/Y _17847_/X VGND VGND VPWR VPWR _17849_/A sky130_fd_sc_hd__or2_4
XFILLER_39_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17779_ _17748_/X _17779_/B _17779_/C VGND VGND VPWR VPWR _17779_/X sky130_fd_sc_hd__and3_4
XANTENNA__22704__B1 _23008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19518_ _21803_/B _19513_/X _11957_/X _19513_/X VGND VGND VPWR VPWR _23720_/D sky130_fd_sc_hd__a2bb2o_4
X_20790_ _20789_/A _20790_/B _20768_/B _13128_/X VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__or4_4
XANTENNA__22180__B2 _14229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19449_ _19448_/Y _19444_/X _19402_/X _19444_/X VGND VGND VPWR VPWR _23744_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_215_0_HCLK clkbuf_8_214_0_HCLK/A VGND VGND VPWR VPWR _25018_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_210_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22460_ _23087_/B VGND VGND VPWR VPWR _22460_/X sky130_fd_sc_hd__buf_2
XFILLER_194_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22019__A _21212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21411_ _21408_/A _21411_/B VGND VGND VPWR VPWR _21411_/X sky130_fd_sc_hd__or2_4
X_22391_ _22387_/X _22390_/X _14686_/X VGND VGND VPWR VPWR _22391_/Y sky130_fd_sc_hd__o21ai_4
X_24130_ _23976_/CLK _18874_/Y HRESETn VGND VGND VPWR VPWR pwm_S7 sky130_fd_sc_hd__dfrtp_4
XFILLER_148_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16698__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21342_ _21311_/A VGND VGND VPWR VPWR _22610_/B sky130_fd_sc_hd__buf_2
XFILLER_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12708__C1 _12662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24061_ _24532_/CLK _20899_/X HRESETn VGND VGND VPWR VPWR _24061_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15856__A _15683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21273_ _21273_/A _21273_/B VGND VGND VPWR VPWR _21275_/B sky130_fd_sc_hd__or2_4
XANTENNA__21577__B _21577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23012_ _16578_/A _22940_/X _22941_/X _23011_/X VGND VGND VPWR VPWR _23013_/C sky130_fd_sc_hd__a211o_4
X_20224_ _21767_/B _20219_/X _19803_/A _20219_/X VGND VGND VPWR VPWR _20224_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_150_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20155_ _20155_/A VGND VGND VPWR VPWR _20155_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22689__A _16284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _20093_/A VGND VGND VPWR VPWR _20086_/X sky130_fd_sc_hd__buf_2
X_24963_ _23991_/CLK _15473_/X HRESETn VGND VGND VPWR VPWR _24963_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_58_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21746__A1 _21565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23914_ _23913_/CLK _23914_/D VGND VGND VPWR VPWR _18965_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24894_ _25062_/CLK _15698_/Y HRESETn VGND VGND VPWR VPWR _24894_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18611__B2 _18737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22201__B _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23845_ _24100_/CLK _23845_/D VGND VGND VPWR VPWR _23845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_25_0_HCLK clkbuf_5_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ HWDATA[20] VGND VGND VPWR VPWR _11790_/X sky130_fd_sc_hd__buf_2
X_23776_ _23850_/CLK _19358_/X VGND VGND VPWR VPWR _18128_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_150_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ scl_oen_o_S4 _20988_/B VGND VGND VPWR VPWR _20988_/X sky130_fd_sc_hd__and2_4
XFILLER_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25515_ _23555_/CLK _25515_/D HRESETn VGND VGND VPWR VPWR _19990_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_213_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22727_ _24874_/Q _22725_/X _21121_/A _22726_/X VGND VGND VPWR VPWR _22728_/C sky130_fd_sc_hd__a211o_4
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24782__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _13428_/A _13460_/B VGND VGND VPWR VPWR _13460_/X sky130_fd_sc_hd__or2_4
X_25446_ _25443_/CLK _12495_/Y HRESETn VGND VGND VPWR VPWR _25446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22658_ _12941_/A _22678_/B _22657_/X VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__o21a_4
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12411_ _12403_/A VGND VGND VPWR VPWR _12411_/X sky130_fd_sc_hd__buf_2
XANTENNA__24711__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21609_ _21121_/X _21604_/Y _21605_/X _21608_/X VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__o22a_4
X_13391_ _13391_/A _13387_/X _13391_/C VGND VGND VPWR VPWR _13391_/X sky130_fd_sc_hd__or3_4
X_25377_ _25380_/CLK _25377_/D HRESETn VGND VGND VPWR VPWR _25377_/Q sky130_fd_sc_hd__dfrtp_4
X_22589_ _16434_/A _22589_/B VGND VGND VPWR VPWR _22592_/B sky130_fd_sc_hd__or2_4
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ _15091_/X _15103_/X _15116_/X _15130_/D VGND VGND VPWR VPWR _15172_/A sky130_fd_sc_hd__or4_4
XFILLER_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12342_ _12342_/A VGND VGND VPWR VPWR _12342_/Y sky130_fd_sc_hd__inv_2
X_24328_ _23654_/CLK _24328_/D HRESETn VGND VGND VPWR VPWR _24328_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15061_ _24471_/Q VGND VGND VPWR VPWR _15061_/Y sky130_fd_sc_hd__inv_2
X_12273_ _12290_/A VGND VGND VPWR VPWR _12273_/X sky130_fd_sc_hd__buf_2
X_24259_ _23494_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _22005_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14012_ _14012_/A _14032_/B _14042_/B _14033_/A VGND VGND VPWR VPWR _14022_/A sky130_fd_sc_hd__or4_4
XFILLER_181_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18820_ _18689_/C _18791_/B VGND VGND VPWR VPWR _18824_/B sky130_fd_sc_hd__or2_4
XANTENNA__17981__A _18097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13286__A _13228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18751_ _18694_/Y _18772_/A _18772_/B VGND VGND VPWR VPWR _18751_/X sky130_fd_sc_hd__or3_4
X_15963_ HWDATA[21] VGND VGND VPWR VPWR _15963_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_214_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16597__A _16618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21737__B2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17702_ _17700_/Y _17702_/B _17702_/C VGND VGND VPWR VPWR _24299_/D sky130_fd_sc_hd__and3_4
XFILLER_208_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14914_ _14914_/A VGND VGND VPWR VPWR _14914_/Y sky130_fd_sc_hd__inv_2
X_15894_ _15713_/X VGND VGND VPWR VPWR _15894_/X sky130_fd_sc_hd__buf_2
X_18682_ _18682_/A VGND VGND VPWR VPWR _18683_/B sky130_fd_sc_hd__buf_2
XFILLER_209_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17633_ _17632_/X VGND VGND VPWR VPWR _24318_/D sky130_fd_sc_hd__inv_2
XFILLER_208_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14845_ _14819_/X _14843_/X _25203_/Q _14844_/X VGND VGND VPWR VPWR _14845_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_224_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14776_ _14779_/A _14781_/A _14776_/C VGND VGND VPWR VPWR _14776_/X sky130_fd_sc_hd__or3_4
X_17564_ _17609_/B VGND VGND VPWR VPWR _17691_/A sky130_fd_sc_hd__buf_2
X_11988_ _11710_/B _11981_/X _11987_/Y VGND VGND VPWR VPWR _11988_/X sky130_fd_sc_hd__a21o_4
XFILLER_189_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19303_ _19299_/Y _19302_/X _19169_/X _19302_/X VGND VGND VPWR VPWR _23796_/D sky130_fd_sc_hd__a2bb2o_4
X_13727_ _11676_/Y _13695_/X VGND VGND VPWR VPWR _13727_/Y sky130_fd_sc_hd__nand2_4
X_16515_ _24565_/Q VGND VGND VPWR VPWR _16515_/Y sky130_fd_sc_hd__inv_2
X_17495_ _17465_/X _17494_/Y _17467_/Y _17494_/A VGND VGND VPWR VPWR _17499_/C sky130_fd_sc_hd__o22a_4
XFILLER_220_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19234_ _20079_/A _20256_/D _20079_/C _18905_/D VGND VGND VPWR VPWR _19234_/X sky130_fd_sc_hd__or4_4
X_13658_ _24064_/Q _20915_/B _24063_/Q _13658_/D VGND VGND VPWR VPWR _13658_/X sky130_fd_sc_hd__or4_4
X_16446_ _16390_/A VGND VGND VPWR VPWR _16446_/X sky130_fd_sc_hd__buf_2
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14564__B _13599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12609_ _12609_/A _12609_/B VGND VGND VPWR VPWR _12609_/X sky130_fd_sc_hd__or2_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16377_ _24616_/Q VGND VGND VPWR VPWR _16377_/Y sky130_fd_sc_hd__inv_2
X_19165_ _23844_/Q VGND VGND VPWR VPWR _19165_/Y sky130_fd_sc_hd__inv_2
X_13589_ _25270_/Q VGND VGND VPWR VPWR _13589_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_45_0_HCLK clkbuf_7_22_0_HCLK/X VGND VGND VPWR VPWR _23493_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_191_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15328_ _15327_/X VGND VGND VPWR VPWR _25011_/D sky130_fd_sc_hd__inv_2
X_18116_ _18227_/A _18112_/X _18115_/X VGND VGND VPWR VPWR _18116_/X sky130_fd_sc_hd__or3_4
XFILLER_118_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19096_ _19095_/Y _19090_/X _18999_/X _19090_/A VGND VGND VPWR VPWR _19096_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15676__A _15676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15259_ _15259_/A _15276_/A _15275_/A _15281_/A VGND VGND VPWR VPWR _15259_/X sky130_fd_sc_hd__or4_4
X_18047_ _18158_/A _18985_/A VGND VGND VPWR VPWR _18048_/C sky130_fd_sc_hd__or2_4
XFILLER_117_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19618__B1 _19454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19148__A _19148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20185__A2_N _20184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18841__A1 _16506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19998_ _22047_/B _19989_/X _19996_/X _19997_/X VGND VGND VPWR VPWR _23554_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16852__B1 _16530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18949_ _18949_/A VGND VGND VPWR VPWR _18949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22302__A _22302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21938_/A _21960_/B VGND VGND VPWR VPWR _21961_/C sky130_fd_sc_hd__or2_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16300__A _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20911_ _20906_/Y _20911_/B _20911_/C VGND VGND VPWR VPWR _20911_/X sky130_fd_sc_hd__and3_4
X_21891_ _12828_/X _21890_/X _24267_/Q _21440_/X VGND VGND VPWR VPWR _21891_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_215_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23630_ _23631_/CLK _23630_/D VGND VGND VPWR VPWR _13435_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _20842_/A VGND VGND VPWR VPWR _20842_/X sky130_fd_sc_hd__buf_2
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20123__A2_N _20118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _23513_/CLK _19975_/X VGND VGND VPWR VPWR _23561_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773_ _20776_/A _20768_/X _20772_/X VGND VGND VPWR VPWR _20773_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18227__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25300_ _24406_/CLK _13710_/Y HRESETn VGND VGND VPWR VPWR _25300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22512_ _14943_/Y _22460_/X _21591_/X _22511_/X VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23516_/CLK _20173_/X VGND VGND VPWR VPWR _20169_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23102__B1 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25231_ _25105_/CLK _14102_/X HRESETn VGND VGND VPWR VPWR _14012_/A sky130_fd_sc_hd__dfrtp_4
X_22443_ _22443_/A VGND VGND VPWR VPWR _22446_/A sky130_fd_sc_hd__buf_2
XFILLER_10_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15591__B1 _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25162_ _25491_/CLK _25162_/D HRESETn VGND VGND VPWR VPWR _25162_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21664__B1 _13804_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22374_ _22085_/A _19786_/Y VGND VGND VPWR VPWR _22374_/X sky130_fd_sc_hd__or2_4
XFILLER_164_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24113_ _23954_/CLK _20978_/Y HRESETn VGND VGND VPWR VPWR _24113_/Q sky130_fd_sc_hd__dfrtp_4
X_21325_ _24048_/Q _21320_/X _21323_/X _21324_/X VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__a211o_4
X_25093_ _25093_/CLK _25093_/D HRESETn VGND VGND VPWR VPWR _25093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14490__A _14485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19609__B1 _19560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24044_ _24509_/CLK _24044_/D HRESETn VGND VGND VPWR VPWR _20822_/A sky130_fd_sc_hd__dfrtp_4
X_21256_ _14687_/A VGND VGND VPWR VPWR _21260_/A sky130_fd_sc_hd__buf_2
XANTENNA__25328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20207_ _23478_/Q VGND VGND VPWR VPWR _21411_/B sky130_fd_sc_hd__inv_2
X_21187_ _21182_/A _21187_/B VGND VGND VPWR VPWR _21187_/X sky130_fd_sc_hd__or2_4
X_20138_ _23504_/Q VGND VGND VPWR VPWR _20138_/Y sky130_fd_sc_hd__inv_2
X_12960_ _12959_/X VGND VGND VPWR VPWR _25383_/D sky130_fd_sc_hd__inv_2
X_20069_ _23528_/Q VGND VGND VPWR VPWR _21788_/B sky130_fd_sc_hd__inv_2
X_24946_ _23407_/CLK _15516_/X HRESETn VGND VGND VPWR VPWR _15515_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23027__B _23027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11911_ RsRx_S1 _11910_/X VGND VGND VPWR VPWR _11911_/X sky130_fd_sc_hd__and2_4
XFILLER_245_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12891_ _12908_/A VGND VGND VPWR VPWR _12891_/X sky130_fd_sc_hd__buf_2
X_24877_ _25433_/CLK _15747_/X HRESETn VGND VGND VPWR VPWR _12568_/A sky130_fd_sc_hd__dfrtp_4
X_14630_ _13647_/X _14629_/X VGND VGND VPWR VPWR _14630_/X sky130_fd_sc_hd__or2_4
XFILLER_61_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11842_ _13844_/A VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__buf_2
X_23828_ _23836_/CLK _23828_/D VGND VGND VPWR VPWR _17951_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14560_/X VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__buf_2
XANTENNA__25150__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ HWDATA[25] VGND VGND VPWR VPWR _11773_/X sky130_fd_sc_hd__buf_2
X_23759_ _23735_/CLK _23759_/D VGND VGND VPWR VPWR _18143_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13512_ _25318_/Q VGND VGND VPWR VPWR _13512_/Y sky130_fd_sc_hd__inv_2
X_16300_ _24645_/Q VGND VGND VPWR VPWR _16300_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17296_/A VGND VGND VPWR VPWR _17280_/X sky130_fd_sc_hd__buf_2
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A VGND VGND VPWR VPWR _21858_/A sky130_fd_sc_hd__inv_2
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22882__A _22155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16231_ _16231_/A VGND VGND VPWR VPWR _16231_/Y sky130_fd_sc_hd__inv_2
X_13443_ _13443_/A _23853_/Q VGND VGND VPWR VPWR _13444_/C sky130_fd_sc_hd__or2_4
X_25429_ _25433_/CLK _25429_/D HRESETn VGND VGND VPWR VPWR _25429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15582__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_4_0_HCLK clkbuf_7_2_0_HCLK/X VGND VGND VPWR VPWR _23407_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_186_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16162_ _16162_/A VGND VGND VPWR VPWR _16162_/X sky130_fd_sc_hd__buf_2
XFILLER_186_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21498__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13374_ _13332_/X _13370_/X _13373_/X VGND VGND VPWR VPWR _13374_/X sky130_fd_sc_hd__or3_4
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15113_ _24988_/Q VGND VGND VPWR VPWR _15401_/A sky130_fd_sc_hd__inv_2
X_12325_ _25359_/Q _24844_/Q _12323_/Y _12324_/Y VGND VGND VPWR VPWR _12335_/A sky130_fd_sc_hd__o22a_4
X_16093_ _24717_/Q VGND VGND VPWR VPWR _16093_/Y sky130_fd_sc_hd__inv_2
X_15044_ _14935_/X _24470_/Q _14935_/X _24470_/Q VGND VGND VPWR VPWR _15044_/X sky130_fd_sc_hd__a2bb2o_4
X_19921_ _19921_/A VGND VGND VPWR VPWR _19921_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12256_ _12255_/Y _24770_/Q _12293_/A _12202_/Y VGND VGND VPWR VPWR _12256_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12699__A1 _12618_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19852_ _19850_/Y _19851_/X _19807_/X _19851_/X VGND VGND VPWR VPWR _19852_/X sky130_fd_sc_hd__a2bb2o_4
X_12187_ _12287_/A _22608_/A _12287_/A _22608_/A VGND VGND VPWR VPWR _12187_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18803_ _18805_/B VGND VGND VPWR VPWR _18803_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20630__A1 _15482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23218__A _23218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19783_ _19782_/Y _19780_/X _19692_/X _19780_/X VGND VGND VPWR VPWR _23630_/D sky130_fd_sc_hd__a2bb2o_4
X_16995_ _24723_/Q _24380_/Q _16080_/Y _17137_/B VGND VGND VPWR VPWR _16995_/X sky130_fd_sc_hd__o22a_4
XFILLER_228_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18734_ _18701_/A _18743_/A VGND VGND VPWR VPWR _18735_/B sky130_fd_sc_hd__or2_4
XANTENNA__17216__A _24351_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15946_ _15945_/Y VGND VGND VPWR VPWR _15947_/A sky130_fd_sc_hd__buf_2
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18665_ _24153_/Q VGND VGND VPWR VPWR _18733_/A sky130_fd_sc_hd__inv_2
XFILLER_236_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20394__B1 _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15877_ _15880_/A VGND VGND VPWR VPWR _15877_/X sky130_fd_sc_hd__buf_2
XFILLER_237_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17616_ _17569_/B _17616_/B VGND VGND VPWR VPWR _17617_/C sky130_fd_sc_hd__or2_4
X_14828_ _14828_/A _14827_/Y _14806_/Y VGND VGND VPWR VPWR _14829_/B sky130_fd_sc_hd__and3_4
XFILLER_221_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18596_ _18594_/Y _18595_/X _18598_/C VGND VGND VPWR VPWR _24166_/D sky130_fd_sc_hd__and3_4
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24633__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17547_ _17547_/A _17544_/X _17545_/X _17546_/X VGND VGND VPWR VPWR _17561_/B sky130_fd_sc_hd__or4_4
X_14759_ _14692_/B _14753_/X VGND VGND VPWR VPWR _14759_/X sky130_fd_sc_hd__and2_4
XFILLER_205_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13820__B1 _13819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17478_ _24213_/Q _17478_/B VGND VGND VPWR VPWR _18905_/D sky130_fd_sc_hd__or2_4
X_19217_ _19225_/A VGND VGND VPWR VPWR _19217_/X sky130_fd_sc_hd__buf_2
X_16429_ _16427_/Y _16423_/X _16241_/X _16428_/X VGND VGND VPWR VPWR _24599_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15573__B1 _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16790__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19148_ _19148_/A VGND VGND VPWR VPWR _19148_/X sky130_fd_sc_hd__buf_2
XFILLER_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19079_ _13213_/B VGND VGND VPWR VPWR _19079_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21110_ _21047_/X _21108_/X _21882_/A _21109_/X VGND VGND VPWR VPWR _21111_/C sky130_fd_sc_hd__a211o_4
XFILLER_145_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22090_ _22090_/A _20107_/Y VGND VGND VPWR VPWR _22091_/C sky130_fd_sc_hd__or2_4
XANTENNA__25421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21041_ _21040_/Y VGND VGND VPWR VPWR _22533_/A sky130_fd_sc_hd__buf_2
XANTENNA__21855__B _21855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24800_ _24781_/CLK _24800_/D HRESETn VGND VGND VPWR VPWR _22564_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22992_ _22991_/X VGND VGND VPWR VPWR _22992_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22967__A _24605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24731_ _24735_/CLK _24731_/D HRESETn VGND VGND VPWR VPWR _24731_/Q sky130_fd_sc_hd__dfrtp_4
X_21943_ _22027_/A VGND VGND VPWR VPWR _21948_/A sky130_fd_sc_hd__buf_2
XFILLER_55_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_7_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19341__A _19048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24662_ _24169_/CLK _16255_/X HRESETn VGND VGND VPWR VPWR _22557_/A sky130_fd_sc_hd__dfrtp_4
X_21874_ _21874_/A VGND VGND VPWR VPWR _23274_/B sky130_fd_sc_hd__buf_2
XFILLER_55_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23615_/CLK _19835_/X VGND VGND VPWR VPWR _23613_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _24045_/Q VGND VGND VPWR VPWR _20825_/Y sky130_fd_sc_hd__inv_2
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24593_ _24989_/CLK _16440_/X HRESETn VGND VGND VPWR VPWR _24593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14485__A _14485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _23560_/CLK _20027_/X VGND VGND VPWR VPWR _23544_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _13142_/D VGND VGND VPWR VPWR _20756_/Y sky130_fd_sc_hd__inv_2
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17189__A2_N _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20077__A2_N _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23475_/CLK _20217_/X VGND VGND VPWR VPWR _20216_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_195_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20687_ _20681_/A _20684_/Y _20685_/Y _20684_/A _20686_/X VGND VGND VPWR VPWR _20687_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25214_ _25212_/CLK _14211_/X HRESETn VGND VGND VPWR VPWR _20511_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22426_ _22296_/X _22424_/X _22298_/X _22425_/X VGND VGND VPWR VPWR _22427_/B sky130_fd_sc_hd__o22a_4
XFILLER_108_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25145_ _25145_/CLK _14436_/X HRESETn VGND VGND VPWR VPWR _25145_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_108_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21111__A _21058_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22357_ _21947_/A _22357_/B VGND VGND VPWR VPWR _22357_/X sky130_fd_sc_hd__or2_4
XFILLER_163_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_91_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _24883_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16205__A _23250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12110_ _12110_/A VGND VGND VPWR VPWR _12123_/A sky130_fd_sc_hd__inv_2
X_21308_ _21320_/A _21307_/X _21308_/C VGND VGND VPWR VPWR _21308_/X sky130_fd_sc_hd__and3_4
XFILLER_123_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13090_ _13004_/B _13089_/X VGND VGND VPWR VPWR _13091_/B sky130_fd_sc_hd__or2_4
X_25076_ _25077_/CLK _25076_/D HRESETn VGND VGND VPWR VPWR _25076_/Q sky130_fd_sc_hd__dfrtp_4
X_22288_ _23093_/A VGND VGND VPWR VPWR _22836_/A sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12041_ _12040_/Y _12038_/X _25498_/Q _12038_/X VGND VGND VPWR VPWR _25499_/D sky130_fd_sc_hd__a2bb2o_4
X_24027_ _24495_/CLK _20751_/X HRESETn VGND VGND VPWR VPWR _13141_/A sky130_fd_sc_hd__dfrtp_4
X_21239_ _21227_/Y _21121_/X _21229_/X _21238_/X VGND VGND VPWR VPWR _21290_/C sky130_fd_sc_hd__a211o_4
XFILLER_151_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15800_ _15800_/A _15934_/B VGND VGND VPWR VPWR _15826_/A sky130_fd_sc_hd__or2_4
XFILLER_172_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13992_ _13992_/A VGND VGND VPWR VPWR _14027_/D sky130_fd_sc_hd__buf_2
X_16780_ _16778_/Y _16779_/X _15761_/X _16779_/X VGND VGND VPWR VPWR _24462_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21781__A _22390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _25386_/Q _12942_/Y VGND VGND VPWR VPWR _12943_/X sky130_fd_sc_hd__or2_4
X_15731_ _12536_/Y _15727_/X _11766_/X _15730_/X VGND VGND VPWR VPWR _15731_/X sky130_fd_sc_hd__a2bb2o_4
X_24929_ _24915_/CLK _24929_/D HRESETn VGND VGND VPWR VPWR _23336_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18450_ _16219_/A _18486_/B _16224_/Y _24183_/Q VGND VGND VPWR VPWR _18451_/D sky130_fd_sc_hd__a2bb2o_4
X_12874_ _12846_/X VGND VGND VPWR VPWR _12908_/A sky130_fd_sc_hd__inv_2
X_15662_ _15661_/X VGND VGND VPWR VPWR _15662_/Y sky130_fd_sc_hd__inv_2
XPHY_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17401_/A _17400_/X VGND VGND VPWR VPWR _17402_/B sky130_fd_sc_hd__or2_4
XPHY_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11803_/X VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__buf_2
X_14613_ _14613_/A _14613_/B VGND VGND VPWR VPWR _14613_/Y sky130_fd_sc_hd__nand2_4
XPHY_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _15592_/Y _15590_/X _11783_/X _15590_/X VGND VGND VPWR VPWR _15593_/X sky130_fd_sc_hd__a2bb2o_4
X_18381_ _24202_/Q VGND VGND VPWR VPWR _18381_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21325__C1 _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20679__A1 _14227_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11812__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14543_/A VGND VGND VPWR VPWR _14544_/Y sky130_fd_sc_hd__inv_2
X_17332_ _17315_/X _17332_/B _17332_/C VGND VGND VPWR VPWR _17332_/X sky130_fd_sc_hd__and3_4
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11754_/Y _11751_/X _11755_/X _11751_/X VGND VGND VPWR VPWR _11756_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _14468_/A VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__buf_2
X_17263_ _17331_/A _17330_/A _17263_/C _17262_/Y VGND VGND VPWR VPWR _17318_/A sky130_fd_sc_hd__or4_4
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11685_/A _24236_/Q _11685_/Y _11686_/Y VGND VGND VPWR VPWR _11687_/X sky130_fd_sc_hd__o22a_4
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19002_ _19166_/A _19166_/B _25079_/Q _19346_/B VGND VGND VPWR VPWR _19002_/X sky130_fd_sc_hd__or4_4
XFILLER_186_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13426_ _13282_/A _19713_/A VGND VGND VPWR VPWR _13426_/X sky130_fd_sc_hd__or2_4
X_16214_ _16214_/A VGND VGND VPWR VPWR _16214_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16951__A2_N _24289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17194_ _24625_/Q _17193_/A _16354_/Y _17193_/Y VGND VGND VPWR VPWR _17200_/B sky130_fd_sc_hd__o22a_4
XFILLER_139_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22825__C1 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16145_ _22649_/A VGND VGND VPWR VPWR _16145_/Y sky130_fd_sc_hd__inv_2
X_13357_ _13421_/A _13357_/B VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__or2_4
XFILLER_6_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22840__A2 _21456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _25365_/Q VGND VGND VPWR VPWR _12308_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16076_ _16004_/X VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__buf_2
XFILLER_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_119_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _25410_/CLK sky130_fd_sc_hd__clkbuf_1
X_13288_ _13245_/X _13288_/B VGND VGND VPWR VPWR _13289_/C sky130_fd_sc_hd__or2_4
XFILLER_170_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15027_ _25043_/Q _15026_/A _14986_/Y _15026_/Y VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__o22a_4
X_19904_ _19904_/A VGND VGND VPWR VPWR _19904_/Y sky130_fd_sc_hd__inv_2
X_12239_ _12255_/A _12237_/Y _12238_/Y _22159_/A VGND VGND VPWR VPWR _12239_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16807__B1 _16385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19835_ _19834_/Y _19829_/X _19761_/X _19816_/A VGND VGND VPWR VPWR _19835_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24885__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19766_ _19765_/Y VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__buf_2
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16978_ _24742_/Q _17105_/A _24748_/Q _17075_/C VGND VGND VPWR VPWR _16980_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22787__A _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21159__A2 _21353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18717_ _18717_/A _18717_/B VGND VGND VPWR VPWR _18720_/B sky130_fd_sc_hd__or2_4
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24814__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15929_ _15686_/X _15928_/Y _15693_/A _15928_/Y VGND VGND VPWR VPWR _24789_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22002__D _22002_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19697_ _18334_/X _20256_/D _19119_/C VGND VGND VPWR VPWR _19698_/A sky130_fd_sc_hd__or3_4
XFILLER_25_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18648_ _18648_/A VGND VGND VPWR VPWR _18809_/A sky130_fd_sc_hd__buf_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18980__B1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18579_ _18556_/X _18573_/B _18578_/Y VGND VGND VPWR VPWR _24172_/D sky130_fd_sc_hd__and3_4
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20610_ _20610_/A _20609_/B VGND VGND VPWR VPWR _20610_/Y sky130_fd_sc_hd__nand2_4
XFILLER_221_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21590_ _14946_/Y _21588_/X _21591_/A _21589_/X VGND VGND VPWR VPWR _21590_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20541_ _20486_/Y _20540_/X _20487_/B VGND VGND VPWR VPWR _20541_/X sky130_fd_sc_hd__o21a_4
XFILLER_138_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15546__B1 HADDR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23260_ _16201_/A _15681_/X VGND VGND VPWR VPWR _23260_/X sky130_fd_sc_hd__or2_4
X_20472_ _20444_/A _20457_/X _20460_/A VGND VGND VPWR VPWR _20473_/B sky130_fd_sc_hd__and3_4
XFILLER_193_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17766__D _16950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22211_ _14765_/X VGND VGND VPWR VPWR _22227_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_180_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22292__B1 _24727_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23191_ _24477_/Q _23016_/X _23190_/X VGND VGND VPWR VPWR _23191_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_78_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22142_ _24489_/Q _22854_/B VGND VGND VPWR VPWR _22145_/B sky130_fd_sc_hd__or2_4
XFILLER_134_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22044__B1 _21697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22073_ _21271_/A VGND VGND VPWR VPWR _22095_/A sky130_fd_sc_hd__buf_2
XFILLER_0_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21024_ _21056_/A _21024_/B VGND VGND VPWR VPWR _21024_/X sky130_fd_sc_hd__and2_4
XFILLER_113_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14285__B1 _13819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22697__A _22535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14199__B _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24555__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22975_ _16125_/Y _22531_/B _15870_/B _11789_/Y _22864_/X VGND VGND VPWR VPWR _22975_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_228_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17223__B1 _24638_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21926_ _22373_/A _21926_/B _21925_/X VGND VGND VPWR VPWR _21926_/X sky130_fd_sc_hd__and3_4
X_24714_ _24697_/CLK _16107_/X HRESETn VGND VGND VPWR VPWR _23237_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24645_ _24639_/CLK _24645_/D HRESETn VGND VGND VPWR VPWR _24645_/Q sky130_fd_sc_hd__dfrtp_4
X_21857_ _16460_/A _21857_/B _21857_/C VGND VGND VPWR VPWR _21880_/A sky130_fd_sc_hd__and3_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _13127_/B VGND VGND VPWR VPWR _20808_/Y sky130_fd_sc_hd__inv_2
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12590_/A VGND VGND VPWR VPWR _12590_/Y sky130_fd_sc_hd__inv_2
X_24576_ _24592_/CLK _24576_/D HRESETn VGND VGND VPWR VPWR _24576_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21788_ _21783_/A _21788_/B VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__or2_4
XFILLER_169_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23527_ _23494_/CLK _20073_/X VGND VGND VPWR VPWR _20071_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ _20788_/A VGND VGND VPWR VPWR _20739_/X sky130_fd_sc_hd__buf_2
XFILLER_211_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14260_/A _14254_/B _15437_/A _14260_/D VGND VGND VPWR VPWR _14260_/X sky130_fd_sc_hd__or4_4
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23458_ _23454_/CLK _23458_/D VGND VGND VPWR VPWR _13275_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13211_ _13211_/A VGND VGND VPWR VPWR _13454_/A sky130_fd_sc_hd__buf_2
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22409_ _22402_/Y _22407_/X _22408_/X _24238_/Q _13828_/D VGND VGND VPWR VPWR _22409_/X
+ sky130_fd_sc_hd__a32o_4
X_14191_ _25135_/Q VGND VGND VPWR VPWR _14191_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14760__A1 _14758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23389_ _23913_/CLK _20435_/X VGND VGND VPWR VPWR _13385_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22822__A2 _22541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13142_ _20752_/A _13141_/X _13142_/C _13142_/D VGND VGND VPWR VPWR _13143_/C sky130_fd_sc_hd__or4_4
X_25128_ _25154_/CLK _25128_/D HRESETn VGND VGND VPWR VPWR _25128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20680__A _20680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13073_ _13069_/A _13066_/X _13072_/Y VGND VGND VPWR VPWR _13073_/X sky130_fd_sc_hd__and3_4
X_17950_ _17950_/A _23836_/Q VGND VGND VPWR VPWR _17950_/X sky130_fd_sc_hd__or2_4
X_25059_ _23385_/CLK _25059_/D HRESETn VGND VGND VPWR VPWR _14812_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__19246__A _19131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ _24108_/Q _12003_/X VGND VGND VPWR VPWR _12024_/X sky130_fd_sc_hd__and2_4
X_16901_ _22199_/A VGND VGND VPWR VPWR _16901_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22586__B2 _22585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17881_ _17881_/A _17877_/X _17880_/Y VGND VGND VPWR VPWR _24269_/D sky130_fd_sc_hd__and3_4
X_19620_ _19761_/A VGND VGND VPWR VPWR _19620_/X sky130_fd_sc_hd__buf_2
X_16832_ _24435_/Q VGND VGND VPWR VPWR _16832_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14276__B1 _13806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _19551_/A VGND VGND VPWR VPWR _19565_/A sky130_fd_sc_hd__buf_2
X_16763_ _16761_/Y _16758_/X _16414_/X _16762_/X VGND VGND VPWR VPWR _16763_/X sky130_fd_sc_hd__a2bb2o_4
X_13975_ _13976_/A _13975_/B VGND VGND VPWR VPWR _13975_/X sky130_fd_sc_hd__and2_4
XANTENNA__22400__A _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18502_ _18492_/A _18500_/X _18502_/C VGND VGND VPWR VPWR _24192_/D sky130_fd_sc_hd__and3_4
XFILLER_234_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ _15713_/X VGND VGND VPWR VPWR _15714_/X sky130_fd_sc_hd__buf_2
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12926_ _12773_/Y _12926_/B VGND VGND VPWR VPWR _12926_/Y sky130_fd_sc_hd__nand2_4
X_19482_ _18282_/X _19480_/X _19481_/X VGND VGND VPWR VPWR _19483_/A sky130_fd_sc_hd__or3_4
X_16694_ _24498_/Q VGND VGND VPWR VPWR _16694_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18962__B1 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18433_ _24164_/Q VGND VGND VPWR VPWR _18433_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15645_ _15645_/A VGND VGND VPWR VPWR _15645_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15776__B1 _24864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12857_ _12857_/A VGND VGND VPWR VPWR _12857_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11808_ HWDATA[15] VGND VGND VPWR VPWR _16238_/A sky130_fd_sc_hd__buf_2
X_18364_ _24206_/Q _17492_/X _18363_/X VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__a21o_4
X_12788_ _22913_/A VGND VGND VPWR VPWR _12788_/Y sky130_fd_sc_hd__inv_2
X_15576_ _24926_/Q VGND VGND VPWR VPWR _23245_/A sky130_fd_sc_hd__inv_2
XANTENNA__17517__A1 _25544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17353_/A VGND VGND VPWR VPWR _17315_/X sky130_fd_sc_hd__buf_2
X_11739_ _11739_/A _11739_/B _11737_/X _11738_/X VGND VGND VPWR VPWR _11740_/D sky130_fd_sc_hd__or4_4
X_14527_ _14524_/A _14525_/X _25126_/Q _14526_/X VGND VGND VPWR VPWR _14527_/X sky130_fd_sc_hd__o22a_4
X_18295_ _18283_/X _18294_/X _18283_/X _18294_/X VGND VGND VPWR VPWR _18295_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17246_ _17310_/A VGND VGND VPWR VPWR _17266_/A sky130_fd_sc_hd__inv_2
X_14458_ _14178_/Y _14457_/X _14404_/X _14457_/X VGND VGND VPWR VPWR _25137_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ _13207_/X _13408_/X _25333_/Q _13267_/X VGND VGND VPWR VPWR _13409_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14389_ _13985_/X _14389_/B VGND VGND VPWR VPWR _14389_/X sky130_fd_sc_hd__or2_4
X_17177_ _17177_/A VGND VGND VPWR VPWR _17178_/A sky130_fd_sc_hd__inv_2
XFILLER_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16128_ _16103_/X VGND VGND VPWR VPWR _16128_/X sky130_fd_sc_hd__buf_2
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16059_ _16058_/Y _16056_/X _15905_/X _16056_/X VGND VGND VPWR VPWR _24731_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19818_ _19814_/Y _19816_/X _19817_/X _19816_/X VGND VGND VPWR VPWR _19818_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17453__B1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11717__A _13782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19749_ _19747_/Y _19743_/X _19659_/X _19748_/X VGND VGND VPWR VPWR _23642_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22760_ _24632_/Q _22610_/B VGND VGND VPWR VPWR _22760_/X sky130_fd_sc_hd__or2_4
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18953__B1 _16861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20355__A3 _15993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14217__A1_N _20525_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _21711_/A _21710_/X VGND VGND VPWR VPWR _21711_/X sky130_fd_sc_hd__and2_4
X_22691_ _11706_/Y _21968_/A _13578_/Y _22523_/A VGND VGND VPWR VPWR _22691_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _24430_/CLK _16847_/X HRESETn VGND VGND VPWR VPWR _16845_/A sky130_fd_sc_hd__dfrtp_4
X_21642_ _22387_/A _21639_/X _21641_/X VGND VGND VPWR VPWR _21642_/X sky130_fd_sc_hd__and3_4
XFILLER_240_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17508__B2 _24312_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24361_ _24346_/CLK _24361_/D HRESETn VGND VGND VPWR VPWR _17340_/A sky130_fd_sc_hd__dfrtp_4
X_21573_ _21566_/Y _21567_/Y _21570_/Y _21572_/Y VGND VGND VPWR VPWR _21573_/X sky130_fd_sc_hd__or4_4
XFILLER_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23312_ _23253_/A _23309_/X _23312_/C VGND VGND VPWR VPWR _23317_/C sky130_fd_sc_hd__and3_4
XFILLER_138_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20524_ _20524_/A _14291_/X _20684_/A VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__and3_4
X_24292_ _24272_/CLK _17789_/X HRESETn VGND VGND VPWR VPWR _17787_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22980__A _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ _23241_/X _23242_/X _22150_/A VGND VGND VPWR VPWR _23243_/X sky130_fd_sc_hd__or3_4
XFILLER_192_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20455_ _20469_/A _20455_/B _20455_/C _20454_/X VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__or4_4
XFILLER_181_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21596__A _21596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23174_ _12299_/A _22998_/X _24289_/Q _22924_/X VGND VGND VPWR VPWR _23174_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20386_ _20385_/Y VGND VGND VPWR VPWR _20386_/X sky130_fd_sc_hd__buf_2
X_22125_ _13514_/Y _12107_/A _12042_/Y _21580_/X VGND VGND VPWR VPWR _22125_/X sky130_fd_sc_hd__o22a_4
XFILLER_134_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_102_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _23386_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24736__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_165_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23916_/CLK sky130_fd_sc_hd__clkbuf_1
X_22056_ _22056_/A _19619_/Y _22055_/X VGND VGND VPWR VPWR _22056_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_8_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21007_ _14832_/A _21006_/X _14804_/Y VGND VGND VPWR VPWR _24006_/D sky130_fd_sc_hd__o21a_4
XFILLER_248_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17444__B1 _16726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13760_ _13759_/Y _13754_/X VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__or2_4
X_22958_ _16322_/A _23027_/B _22830_/C VGND VGND VPWR VPWR _22958_/X sky130_fd_sc_hd__and3_4
XFILLER_244_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12711_ _12740_/A _12742_/A _12737_/A _12737_/B VGND VGND VPWR VPWR _12712_/B sky130_fd_sc_hd__or4_4
X_21909_ _22093_/A _21909_/B VGND VGND VPWR VPWR _21909_/X sky130_fd_sc_hd__or2_4
X_13691_ _13691_/A _13690_/X VGND VGND VPWR VPWR _13691_/X sky130_fd_sc_hd__or2_4
XFILLER_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22889_ _22887_/X _22888_/X _22510_/C VGND VGND VPWR VPWR _22889_/X sky130_fd_sc_hd__or3_4
XFILLER_204_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12642_ _12642_/A _12642_/B _12702_/A _12642_/D VGND VGND VPWR VPWR _12642_/X sky130_fd_sc_hd__or4_4
X_15430_ _15423_/B VGND VGND VPWR VPWR _15430_/Y sky130_fd_sc_hd__inv_2
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24628_ _24625_/CLK _16347_/X HRESETn VGND VGND VPWR VPWR _24628_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15306_/X _15360_/X VGND VGND VPWR VPWR _15361_/X sky130_fd_sc_hd__or2_4
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _25407_/Q _12571_/Y _25411_/Q _12572_/Y VGND VGND VPWR VPWR _12578_/B sky130_fd_sc_hd__a2bb2o_4
X_24559_ _24556_/CLK _24559_/D HRESETn VGND VGND VPWR VPWR _16529_/A sky130_fd_sc_hd__dfrtp_4
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ _17032_/Y _17086_/B VGND VGND VPWR VPWR _17101_/B sky130_fd_sc_hd__or2_4
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14312_ _14303_/A _14303_/B _13649_/X _14311_/X VGND VGND VPWR VPWR _14313_/A sky130_fd_sc_hd__a211o_4
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _15292_/A _15256_/X VGND VGND VPWR VPWR _15292_/Y sky130_fd_sc_hd__nand2_4
X_18080_ _18209_/A _18080_/B VGND VGND VPWR VPWR _18082_/B sky130_fd_sc_hd__or2_4
XFILLER_183_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22890__A _16684_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21059__A1 _24860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14242_/Y _14238_/X _13809_/X _14238_/X VGND VGND VPWR VPWR _14243_/X sky130_fd_sc_hd__a2bb2o_4
X_17031_ _24408_/Q VGND VGND VPWR VPWR _17060_/A sky130_fd_sc_hd__inv_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15930__B1 _15686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14174_ _14174_/A _14174_/B _14190_/A _14131_/X VGND VGND VPWR VPWR _14174_/X sky130_fd_sc_hd__or4_4
XANTENNA__19672__B2 _19652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_61_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13125_ _13088_/A _13026_/D _13019_/A _13123_/B VGND VGND VPWR VPWR _13126_/A sky130_fd_sc_hd__a211o_4
X_18982_ _18981_/Y _14674_/X _17427_/X _14674_/X VGND VGND VPWR VPWR _23908_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22559__A1 _16522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _25361_/Q _13055_/Y VGND VGND VPWR VPWR _13056_/X sky130_fd_sc_hd__or2_4
X_17933_ _17929_/Y _17924_/B VGND VGND VPWR VPWR _17933_/X sky130_fd_sc_hd__or2_4
XFILLER_140_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23220__A2 _22485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12640__B _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12007_ _12000_/X VGND VGND VPWR VPWR _12007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17435__B1 _17433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17864_ _17864_/A _17864_/B VGND VGND VPWR VPWR _17865_/C sky130_fd_sc_hd__or2_4
XANTENNA__19704__A _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14249__B1 _14248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19603_ _21981_/B VGND VGND VPWR VPWR _19603_/Y sky130_fd_sc_hd__inv_2
X_16815_ _24445_/Q VGND VGND VPWR VPWR _16815_/Y sky130_fd_sc_hd__inv_2
X_17795_ _16910_/A _17800_/B VGND VGND VPWR VPWR _17797_/B sky130_fd_sc_hd__or2_4
XANTENNA__15997__B1 _15848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19534_ _19528_/Y VGND VGND VPWR VPWR _19534_/X sky130_fd_sc_hd__buf_2
XFILLER_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16746_ _16745_/Y _16743_/X _16393_/X _16743_/X VGND VGND VPWR VPWR _24479_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13958_ _13958_/A _13941_/Y _13933_/X _13957_/Y VGND VGND VPWR VPWR _13958_/X sky130_fd_sc_hd__and4_4
XFILLER_47_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22731__A1 _16140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22731__B2 _22289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12909_ _12908_/X VGND VGND VPWR VPWR _25395_/D sky130_fd_sc_hd__inv_2
X_19465_ _18046_/B VGND VGND VPWR VPWR _19465_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16677_ _16677_/A VGND VGND VPWR VPWR _16677_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13889_ _25250_/Q _13869_/X _21160_/A _13864_/X VGND VGND VPWR VPWR _13889_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18416_ _24187_/Q VGND VGND VPWR VPWR _18517_/A sky130_fd_sc_hd__inv_2
XFILLER_50_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15628_ _24905_/Q VGND VGND VPWR VPWR _15628_/Y sky130_fd_sc_hd__inv_2
X_19396_ _23762_/Q VGND VGND VPWR VPWR _19396_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14421__B1 _14420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ _18347_/A _18347_/B VGND VGND VPWR VPWR _18347_/X sky130_fd_sc_hd__or2_4
XANTENNA__15679__A _21170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ _14385_/A _16378_/B _16190_/C _15559_/D VGND VGND VPWR VPWR _21122_/A sky130_fd_sc_hd__or4_4
XFILLER_159_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18278_ _18277_/X VGND VGND VPWR VPWR _18278_/X sky130_fd_sc_hd__buf_2
XANTENNA__16174__B1 _15848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17229_ _17229_/A VGND VGND VPWR VPWR _17229_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20240_ _20234_/Y VGND VGND VPWR VPWR _20240_/X sky130_fd_sc_hd__buf_2
XFILLER_174_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20171_ _20170_/X VGND VGND VPWR VPWR _20172_/A sky130_fd_sc_hd__inv_2
XFILLER_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14488__B1 _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_238_0_HCLK clkbuf_8_238_0_HCLK/A VGND VGND VPWR VPWR _25105_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23930_ _23514_/CLK _23930_/D VGND VGND VPWR VPWR _23930_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23861_ _23445_/CLK _19117_/X VGND VGND VPWR VPWR _23861_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23136__A _22535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15988__B1 _15629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22040__A _22029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14758__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19179__B1 _19131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22812_ _22811_/X VGND VGND VPWR VPWR _22813_/A sky130_fd_sc_hd__inv_2
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23792_ _23794_/CLK _19314_/X VGND VGND VPWR VPWR _23792_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22722__A1 _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22743_ _22592_/A _22743_/B _22743_/C VGND VGND VPWR VPWR _22743_/X sky130_fd_sc_hd__and3_4
X_25531_ _25528_/CLK _25531_/D HRESETn VGND VGND VPWR VPWR _25531_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12278__A _25444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22694__B _22694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25462_ _25380_/CLK _12431_/Y HRESETn VGND VGND VPWR VPWR _25462_/Q sky130_fd_sc_hd__dfrtp_4
X_22674_ _15718_/A _22673_/X _22148_/C _11816_/A _22695_/B VGND VGND VPWR VPWR _22674_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23278__A2 _23269_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15755__A3 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24413_ _23799_/CLK _24413_/D HRESETn VGND VGND VPWR VPWR _20119_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_213_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21625_ _21625_/A _21625_/B VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__or2_4
XANTENNA__22486__B1 _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25393_ _25402_/CLK _25393_/D HRESETn VGND VGND VPWR VPWR _25393_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19351__B1 _19305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24344_ _24343_/CLK _24344_/D HRESETn VGND VGND VPWR VPWR _24344_/Q sky130_fd_sc_hd__dfstp_4
X_21556_ _21554_/X _21555_/X _21113_/X VGND VGND VPWR VPWR _21556_/X sky130_fd_sc_hd__or3_4
XFILLER_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16165__B1 _16073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17300__C _17355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24329__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20507_ _14214_/A _20505_/X _20499_/C _20506_/X VGND VGND VPWR VPWR _20508_/B sky130_fd_sc_hd__a22oi_4
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24275_ _24272_/CLK _17854_/Y HRESETn VGND VGND VPWR VPWR _24275_/Q sky130_fd_sc_hd__dfrtp_4
X_21487_ _21679_/A _21487_/B _21487_/C VGND VGND VPWR VPWR _21487_/X sky130_fd_sc_hd__or3_4
X_23226_ _23156_/A _23217_/Y _23221_/X _23226_/D VGND VGND VPWR VPWR _23226_/X sky130_fd_sc_hd__or4_4
XFILLER_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20438_ _20438_/A _20475_/C VGND VGND VPWR VPWR _20438_/X sky130_fd_sc_hd__or2_4
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_48_0_HCLK clkbuf_5_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21461__A1 _22810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23157_ _23132_/X _23135_/X _23142_/Y _23156_/X VGND VGND VPWR VPWR HRDATA[25] sky130_fd_sc_hd__a211o_4
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16735__A2_N _16734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21461__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20369_ _20369_/A VGND VGND VPWR VPWR _20369_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22108_ _22941_/A VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__buf_2
XFILLER_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24570__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23088_ _16571_/A _22411_/X _15676_/X _23087_/X VGND VGND VPWR VPWR _23088_/X sky130_fd_sc_hd__a211o_4
XFILLER_164_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15140__B2 _16427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14930_ _25020_/Q VGND VGND VPWR VPWR _14930_/Y sky130_fd_sc_hd__inv_2
X_22039_ _22028_/A _22039_/B VGND VGND VPWR VPWR _22040_/C sky130_fd_sc_hd__or2_4
XFILLER_88_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22961__A1 _12834_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14861_ _14824_/A _14824_/B _14824_/A _14824_/B VGND VGND VPWR VPWR _14862_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_248_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16600_ _16599_/Y _16597_/X _16245_/X _16597_/X VGND VGND VPWR VPWR _24533_/D sky130_fd_sc_hd__a2bb2o_4
X_13812_ _15486_/A VGND VGND VPWR VPWR _13812_/X sky130_fd_sc_hd__buf_2
XFILLER_235_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17580_ _17666_/A VGND VGND VPWR VPWR _17667_/A sky130_fd_sc_hd__inv_2
X_14792_ _14785_/X VGND VGND VPWR VPWR _14792_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14651__B1 _18069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15994__A3 _15993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16531_ _16529_/Y _16525_/X _16530_/X _16525_/X VGND VGND VPWR VPWR _24559_/D sky130_fd_sc_hd__a2bb2o_4
X_13743_ _25285_/Q VGND VGND VPWR VPWR _13744_/A sky130_fd_sc_hd__inv_2
XANTENNA__12188__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19250_ _19248_/Y _19249_/X _19226_/X _19249_/X VGND VGND VPWR VPWR _23815_/D sky130_fd_sc_hd__a2bb2o_4
X_16462_ _13821_/B _21580_/A _16462_/C _15661_/C VGND VGND VPWR VPWR _16462_/X sky130_fd_sc_hd__or4_4
X_13674_ _13673_/X VGND VGND VPWR VPWR _13674_/X sky130_fd_sc_hd__buf_2
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18201_ _18169_/A _18201_/B _18200_/X VGND VGND VPWR VPWR _18202_/C sky130_fd_sc_hd__and3_4
XFILLER_232_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15413_ _15401_/A _15401_/B VGND VGND VPWR VPWR _15413_/Y sky130_fd_sc_hd__nand2_4
X_12625_ _12713_/A _12590_/Y _12737_/A _12538_/Y VGND VGND VPWR VPWR _12626_/C sky130_fd_sc_hd__or4_4
X_19181_ _19181_/A VGND VGND VPWR VPWR _19181_/X sky130_fd_sc_hd__buf_2
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16393_ HWDATA[28] VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__buf_2
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12916__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19342__B1 _19341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18132_ _18164_/A _23848_/Q VGND VGND VPWR VPWR _18134_/B sky130_fd_sc_hd__or2_4
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12556_ _12644_/A _24889_/Q _12631_/C _12555_/Y VGND VGND VPWR VPWR _12566_/A sky130_fd_sc_hd__o22a_4
X_15344_ _15343_/X VGND VGND VPWR VPWR _25007_/D sky130_fd_sc_hd__inv_2
XFILLER_200_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ _18063_/A _18060_/X _18063_/C VGND VGND VPWR VPWR _18063_/X sky130_fd_sc_hd__and3_4
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12288_/Y _12486_/X _12421_/A _12482_/Y VGND VGND VPWR VPWR _12488_/A sky130_fd_sc_hd__a211o_4
X_15275_ _15275_/A _15281_/A VGND VGND VPWR VPWR _15276_/B sky130_fd_sc_hd__or2_4
XFILLER_8_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15903__B1 _22605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17014_ _24406_/Q VGND VGND VPWR VPWR _17034_/A sky130_fd_sc_hd__inv_2
X_14226_ _14225_/Y _14210_/A _13809_/X _14210_/A VGND VGND VPWR VPWR _14226_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24658__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ _14157_/A VGND VGND VPWR VPWR _14157_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ _13051_/A VGND VGND VPWR VPWR _13121_/C sky130_fd_sc_hd__buf_2
X_14088_ _13999_/C _14074_/X _14087_/X _14013_/B _14085_/X VGND VGND VPWR VPWR _25241_/D
+ sky130_fd_sc_hd__a32o_4
X_18965_ _18965_/A VGND VGND VPWR VPWR _18965_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _12329_/Y _13039_/B VGND VGND VPWR VPWR _13044_/B sky130_fd_sc_hd__or2_4
X_17916_ _17908_/Y _17915_/A _17914_/X _17900_/A _17915_/Y VGND VGND VPWR VPWR _17916_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15962__A _15947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18896_ _18876_/X _18890_/X _23966_/Q _24127_/Q _18893_/X VGND VGND VPWR VPWR _18896_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_121_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17847_ _17609_/B _17761_/X VGND VGND VPWR VPWR _17847_/X sky130_fd_sc_hd__or2_4
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_68_0_HCLK clkbuf_7_34_0_HCLK/X VGND VGND VPWR VPWR _25456_/CLK sky130_fd_sc_hd__clkbuf_1
X_17778_ _23332_/A _17776_/Y VGND VGND VPWR VPWR _17779_/C sky130_fd_sc_hd__nand2_4
XFILLER_208_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22704__A1 _22479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19517_ _23720_/Q VGND VGND VPWR VPWR _21803_/B sky130_fd_sc_hd__inv_2
XFILLER_223_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22704__B2 _22703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16729_ _16729_/A VGND VGND VPWR VPWR _16729_/X sky130_fd_sc_hd__buf_2
XFILLER_222_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19448_ _18118_/B VGND VGND VPWR VPWR _19448_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16813__A1_N _14976_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19379_ _23768_/Q VGND VGND VPWR VPWR _19379_/Y sky130_fd_sc_hd__inv_2
X_21410_ _14688_/X _21410_/B VGND VGND VPWR VPWR _21410_/X sky130_fd_sc_hd__or2_4
X_22390_ _22390_/A _22390_/B _22390_/C VGND VGND VPWR VPWR _22390_/X sky130_fd_sc_hd__and3_4
X_21341_ _21235_/X VGND VGND VPWR VPWR _21341_/X sky130_fd_sc_hd__buf_2
X_24060_ _24532_/CLK _20894_/X HRESETn VGND VGND VPWR VPWR _13672_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21272_ _21638_/A _21272_/B _21272_/C VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__and3_4
XFILLER_163_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23011_ _24573_/Q _22897_/X _22816_/X VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__o21a_4
X_20223_ _20223_/A VGND VGND VPWR VPWR _21767_/B sky130_fd_sc_hd__inv_2
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12561__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20154_ _20153_/Y _20151_/X _20105_/X _20151_/X VGND VGND VPWR VPWR _20154_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15122__B2 _15121_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21593__B _21752_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20085_ _13282_/B VGND VGND VPWR VPWR _20085_/Y sky130_fd_sc_hd__inv_2
X_24962_ _23991_/CLK _15475_/X HRESETn VGND VGND VPWR VPWR _24962_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23913_ _23913_/CLK _23913_/D VGND VGND VPWR VPWR _23913_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_218_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24893_ _25062_/CLK _15706_/X HRESETn VGND VGND VPWR VPWR _24893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20954__B1 _20836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23844_ _23836_/CLK _19170_/X VGND VGND VPWR VPWR _23844_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15976__A3 HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ _23889_/CLK _19361_/X VGND VGND VPWR VPWR _23775_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ _20987_/A VGND VGND VPWR VPWR _20988_/B sky130_fd_sc_hd__inv_2
XFILLER_214_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25514_ _23555_/CLK _11940_/X HRESETn VGND VGND VPWR VPWR _19993_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22726_ _22726_/A _21877_/B _21096_/X VGND VGND VPWR VPWR _22726_/X sky130_fd_sc_hd__and3_4
XANTENNA__16386__B1 _16385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23313__B _23313_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20182__B2 _20177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22657_ _17763_/Y _21457_/X _12439_/B _22447_/A VGND VGND VPWR VPWR _22657_/X sky130_fd_sc_hd__o22a_4
X_25445_ _24765_/CLK _12499_/X HRESETn VGND VGND VPWR VPWR _12218_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12410_ _12398_/A _12410_/B _12409_/X VGND VGND VPWR VPWR _12410_/X sky130_fd_sc_hd__and3_4
X_21608_ _13660_/Y _21606_/X _24017_/Q _21607_/X VGND VGND VPWR VPWR _21608_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _13454_/A _13390_/B _13390_/C VGND VGND VPWR VPWR _13391_/C sky130_fd_sc_hd__and3_4
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22588_ _22548_/X _22556_/Y _22588_/C _22587_/Y VGND VGND VPWR VPWR HRDATA[10] sky130_fd_sc_hd__or4_4
X_25376_ _24792_/CLK _12982_/X HRESETn VGND VGND VPWR VPWR _25376_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21131__B1 _21129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12341_ _25349_/Q _24834_/Q _12339_/Y _12340_/Y VGND VGND VPWR VPWR _12341_/X sky130_fd_sc_hd__o22a_4
X_21539_ _21530_/X _21537_/X _21532_/X _12561_/A _21538_/X VGND VGND VPWR VPWR _21540_/B
+ sky130_fd_sc_hd__a32o_4
X_24327_ _24327_/CLK _24327_/D HRESETn VGND VGND VPWR VPWR _17596_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20672__B _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15060_ _24477_/Q VGND VGND VPWR VPWR _15060_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24751__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12272_ _12272_/A VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__inv_2
X_24258_ _24258_/CLK _17927_/X HRESETn VGND VGND VPWR VPWR _24258_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14011_ _14011_/A _13992_/A _25238_/Q _14011_/D VGND VGND VPWR VPWR _14033_/A sky130_fd_sc_hd__or4_4
XANTENNA__15900__A3 _16245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23209_ _12191_/Y _22998_/X _16910_/A _22501_/X VGND VGND VPWR VPWR _23209_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24189_ _24189_/CLK _24189_/D HRESETn VGND VGND VPWR VPWR _24189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21784__A _22387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16310__B1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12388__A2_N _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18750_ _18699_/A _18699_/B _18733_/C _18700_/A VGND VGND VPWR VPWR _18772_/B sky130_fd_sc_hd__or4_4
XANTENNA__15782__A _19761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19254__A _19139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15962_ _15947_/A VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__buf_2
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_221_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _25011_/CLK sky130_fd_sc_hd__clkbuf_1
X_17701_ _17701_/A _17701_/B VGND VGND VPWR VPWR _17702_/B sky130_fd_sc_hd__or2_4
XFILLER_248_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14913_ _24440_/Q VGND VGND VPWR VPWR _14913_/Y sky130_fd_sc_hd__inv_2
X_18681_ _18681_/A VGND VGND VPWR VPWR _18681_/Y sky130_fd_sc_hd__inv_2
X_15893_ _12801_/Y _15890_/X _11800_/X _15890_/X VGND VGND VPWR VPWR _15893_/X sky130_fd_sc_hd__a2bb2o_4
X_17632_ _17895_/B _17629_/B _17632_/C VGND VGND VPWR VPWR _17632_/X sky130_fd_sc_hd__or3_4
XFILLER_236_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14844_ _14835_/A VGND VGND VPWR VPWR _14844_/X sky130_fd_sc_hd__buf_2
XFILLER_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17563_ _17562_/X VGND VGND VPWR VPWR _17609_/B sky130_fd_sc_hd__buf_2
X_14775_ _13749_/Y _14775_/B VGND VGND VPWR VPWR _14776_/C sky130_fd_sc_hd__and2_4
XFILLER_17_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11987_ _11985_/X VGND VGND VPWR VPWR _11987_/Y sky130_fd_sc_hd__inv_2
X_19302_ _19301_/Y VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__buf_2
XFILLER_17_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19563__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16514_ _16512_/Y _16508_/X _16241_/X _16513_/X VGND VGND VPWR VPWR _24566_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13726_ _13698_/B _13716_/X _13725_/Y _13723_/X _11694_/A VGND VGND VPWR VPWR _13726_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_204_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17494_ _17494_/A VGND VGND VPWR VPWR _17494_/Y sky130_fd_sc_hd__inv_2
X_19233_ _18332_/A VGND VGND VPWR VPWR _20256_/D sky130_fd_sc_hd__buf_2
XFILLER_220_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16445_ _16445_/A VGND VGND VPWR VPWR _16445_/Y sky130_fd_sc_hd__inv_2
X_13657_ _24074_/Q _24073_/Q VGND VGND VPWR VPWR _13675_/C sky130_fd_sc_hd__or2_4
X_12608_ _12608_/A _12608_/B _12608_/C _12608_/D VGND VGND VPWR VPWR _12609_/B sky130_fd_sc_hd__or4_4
X_19164_ _19163_/Y _19159_/X _19139_/X _19159_/A VGND VGND VPWR VPWR _23845_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16129__B1 _15967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24839__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16376_ _16374_/Y _16291_/A _16375_/X _16291_/A VGND VGND VPWR VPWR _24617_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13588_ _25097_/Q VGND VGND VPWR VPWR _14601_/A sky130_fd_sc_hd__inv_2
X_18115_ _17988_/A _18115_/B _18115_/C VGND VGND VPWR VPWR _18115_/X sky130_fd_sc_hd__and3_4
X_15327_ _15324_/X _15321_/B _15327_/C VGND VGND VPWR VPWR _15327_/X sky130_fd_sc_hd__or3_4
XFILLER_157_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15957__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12539_ _12538_/Y _24860_/Q _12538_/Y _24860_/Q VGND VGND VPWR VPWR _12540_/D sky130_fd_sc_hd__a2bb2o_4
X_19095_ _13442_/B VGND VGND VPWR VPWR _19095_/Y sky130_fd_sc_hd__inv_2
XFILLER_219_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17558__A1_N _25553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18046_ _18189_/A _18046_/B VGND VGND VPWR VPWR _18046_/X sky130_fd_sc_hd__or2_4
X_15258_ _15258_/A _15257_/X VGND VGND VPWR VPWR _15281_/A sky130_fd_sc_hd__or2_4
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ _14209_/A VGND VGND VPWR VPWR _14210_/A sky130_fd_sc_hd__buf_2
XFILLER_99_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13477__A _21577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15189_ _15182_/A _15186_/X VGND VGND VPWR VPWR _15190_/C sky130_fd_sc_hd__or2_4
XANTENNA__21694__A _21668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16301__B1 _15950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19997_ _19988_/Y VGND VGND VPWR VPWR _19997_/X sky130_fd_sc_hd__buf_2
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18948_ _18947_/Y _18945_/X _16791_/X _18945_/X VGND VGND VPWR VPWR _23921_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22302__B _21091_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22925__B2 _22924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18879_ _20566_/A _18878_/X VGND VGND VPWR VPWR _20567_/A sky130_fd_sc_hd__or2_4
XFILLER_227_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20910_ _24064_/Q VGND VGND VPWR VPWR _20911_/C sky130_fd_sc_hd__inv_2
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21890_ _21027_/X VGND VGND VPWR VPWR _21890_/X sky130_fd_sc_hd__buf_2
XFILLER_215_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20841_ _20840_/X VGND VGND VPWR VPWR _24048_/D sky130_fd_sc_hd__inv_2
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23560_ _23560_/CLK _19977_/X VGND VGND VPWR VPWR _19976_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_223_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20772_ _20772_/A _20763_/Y _20772_/C VGND VGND VPWR VPWR _20772_/X sky130_fd_sc_hd__and3_4
XANTENNA__20164__B2 _20163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22511_ _15022_/Y _22513_/B VGND VGND VPWR VPWR _22511_/X sky130_fd_sc_hd__and2_4
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23516_/CLK _20175_/X VGND VGND VPWR VPWR _23491_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19306__B1 _19305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22442_ _22442_/A _22442_/B VGND VGND VPWR VPWR _22452_/B sky130_fd_sc_hd__nor2_4
X_25230_ _23395_/CLK _14130_/X HRESETn VGND VGND VPWR VPWR _25230_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19857__B2 _19838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25161_ _25168_/CLK _14378_/X HRESETn VGND VGND VPWR VPWR _25161_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22373_ _22373_/A _22371_/X _22372_/X VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__and3_4
XANTENNA__15867__A _15866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_227_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24112_ _24112_/CLK _14340_/Y HRESETn VGND VGND VPWR VPWR _14359_/A sky130_fd_sc_hd__dfrtp_4
X_21324_ _21064_/X VGND VGND VPWR VPWR _21324_/X sky130_fd_sc_hd__buf_2
XFILLER_136_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25092_ _25309_/CLK _14614_/X HRESETn VGND VGND VPWR VPWR _25092_/Q sky130_fd_sc_hd__dfrtp_4
X_24043_ _24509_/CLK _20820_/X HRESETn VGND VGND VPWR VPWR _20822_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21255_ _21638_/A _21253_/X _21254_/X VGND VGND VPWR VPWR _21255_/X sky130_fd_sc_hd__and3_4
XFILLER_190_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20292__A2_N _20291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20206_ _20204_/Y _20205_/X _20119_/X _20205_/X VGND VGND VPWR VPWR _23479_/D sky130_fd_sc_hd__a2bb2o_4
X_21186_ _21207_/A _19921_/Y VGND VGND VPWR VPWR _21188_/B sky130_fd_sc_hd__or2_4
XFILLER_132_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20137_ _21910_/B _20134_/X _20112_/X _20134_/X VGND VGND VPWR VPWR _23505_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16705__A1_N _16703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22212__B _20104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20068_ _21922_/B _20065_/X _19800_/X _20065_/X VGND VGND VPWR VPWR _20068_/X sky130_fd_sc_hd__a2bb2o_4
X_24945_ _23407_/CLK _24945_/D HRESETn VGND VGND VPWR VPWR _15517_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23027__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11910_ _11910_/A VGND VGND VPWR VPWR _11910_/X sky130_fd_sc_hd__buf_2
XFILLER_161_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12890_ _12906_/A _12890_/B _12889_/X VGND VGND VPWR VPWR _25400_/D sky130_fd_sc_hd__and3_4
X_24876_ _24872_/CLK _24876_/D HRESETn VGND VGND VPWR VPWR _24876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_51_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _24406_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_233_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23324__A _21714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ HWDATA[7] VGND VGND VPWR VPWR _13844_/A sky130_fd_sc_hd__buf_2
X_23827_ _23850_/CLK _23827_/D VGND VGND VPWR VPWR _19214_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17322__A _17322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _25550_/Q VGND VGND VPWR VPWR _11772_/Y sky130_fd_sc_hd__inv_2
X_14560_ HSEL VGND VGND VPWR VPWR _14560_/X sky130_fd_sc_hd__buf_2
XFILLER_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12093__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23758_ _23735_/CLK _23758_/D VGND VGND VPWR VPWR _18175_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _11999_/Y _13507_/X _11842_/X _13510_/X VGND VGND VPWR VPWR _13511_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ _20895_/Y _21605_/X _16694_/Y _22460_/X VGND VGND VPWR VPWR _22709_/X sky130_fd_sc_hd__o22a_4
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14489_/Y _14485_/X _14427_/X _14490_/X VGND VGND VPWR VPWR _14491_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23689_ _24206_/CLK _19609_/X VGND VGND VPWR VPWR _19608_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_198_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16230_ _16229_/Y _16227_/X _15970_/X _16227_/X VGND VGND VPWR VPWR _16230_/X sky130_fd_sc_hd__a2bb2o_4
X_13442_ _13410_/A _13442_/B VGND VGND VPWR VPWR _13444_/B sky130_fd_sc_hd__or2_4
X_25428_ _25433_/CLK _25428_/D HRESETn VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21779__A _22388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13373_ _13469_/A _13373_/B _13373_/C VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__and3_4
X_16161_ _22201_/A VGND VGND VPWR VPWR _16161_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15777__A _11861_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25359_ _25425_/CLK _25359_/D HRESETn VGND VGND VPWR VPWR _25359_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_24_0_HCLK_A clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _25005_/Q _24609_/Q _15347_/A _15111_/Y VGND VGND VPWR VPWR _15112_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12324_ _24844_/Q VGND VGND VPWR VPWR _12324_/Y sky130_fd_sc_hd__inv_2
X_16092_ _11730_/Y _21596_/A _16090_/X _24718_/Q _16091_/X VGND VGND VPWR VPWR _24718_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16531__B1 _16530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12255_ _12255_/A VGND VGND VPWR VPWR _12255_/Y sky130_fd_sc_hd__inv_2
X_15043_ _15079_/A _16754_/A _15079_/A _16754_/A VGND VGND VPWR VPWR _15043_/X sky130_fd_sc_hd__a2bb2o_4
X_19920_ _21495_/B _19917_/X _19646_/X _19917_/X VGND VGND VPWR VPWR _23582_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17992__A _18006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19851_ _19838_/Y VGND VGND VPWR VPWR _19851_/X sky130_fd_sc_hd__buf_2
X_12186_ _25449_/Q VGND VGND VPWR VPWR _12287_/A sky130_fd_sc_hd__inv_2
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_36_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__20091__B1 _19753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18802_ _18799_/B _18799_/C VGND VGND VPWR VPWR _18805_/B sky130_fd_sc_hd__or2_4
X_19782_ _13435_/B VGND VGND VPWR VPWR _19782_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16994_ _24380_/Q VGND VGND VPWR VPWR _17137_/B sky130_fd_sc_hd__inv_2
XANTENNA__13648__A1 _13547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18733_ _18733_/A _18733_/B _18733_/C VGND VGND VPWR VPWR _18743_/A sky130_fd_sc_hd__or3_4
X_15945_ _15939_/X VGND VGND VPWR VPWR _15945_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15929__A1_N _15686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18664_ _16566_/Y _24157_/Q _24540_/Q _18696_/D VGND VGND VPWR VPWR _18664_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15876_ _15875_/Y VGND VGND VPWR VPWR _15880_/A sky130_fd_sc_hd__buf_2
XANTENNA__16598__B1 _16241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17615_ _17512_/A _17615_/B VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__or2_4
X_14827_ _14826_/X VGND VGND VPWR VPWR _14827_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22776__C _22754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23234__A _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18595_ _18595_/A _18598_/A VGND VGND VPWR VPWR _18595_/X sky130_fd_sc_hd__or2_4
XFILLER_205_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12265__A2_N _24757_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17546_ _11807_/Y _17575_/A _11807_/Y _17575_/A VGND VGND VPWR VPWR _17546_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12084__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14758_ _22221_/A VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__buf_2
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13709_ _11682_/Y _13705_/A _13708_/X _13703_/X VGND VGND VPWR VPWR _13710_/A sky130_fd_sc_hd__o22a_4
X_17477_ _17477_/A _17477_/B VGND VGND VPWR VPWR _20079_/D sky130_fd_sc_hd__or2_4
X_14689_ _14688_/X VGND VGND VPWR VPWR _21257_/A sky130_fd_sc_hd__buf_2
XFILLER_177_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22792__B _22662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19216_ _18066_/B VGND VGND VPWR VPWR _19216_/Y sky130_fd_sc_hd__inv_2
X_16428_ _16442_/A VGND VGND VPWR VPWR _16428_/X sky130_fd_sc_hd__buf_2
XANTENNA__21689__A _22029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24673__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19147_ _23851_/Q VGND VGND VPWR VPWR _19147_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24602__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _16352_/A VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__buf_2
XANTENNA__19159__A _19159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19078_ _19074_/Y _19077_/X _19032_/X _19077_/X VGND VGND VPWR VPWR _19078_/X sky130_fd_sc_hd__a2bb2o_4
X_18029_ _18029_/A VGND VGND VPWR VPWR _18029_/X sky130_fd_sc_hd__buf_2
X_21040_ _21032_/X VGND VGND VPWR VPWR _21040_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21855__C _21752_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20082__B1 _19817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22991_ _22788_/X _22989_/X _22497_/X _24742_/Q _22990_/X VGND VGND VPWR VPWR _22991_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24730_ _24735_/CLK _16062_/X HRESETn VGND VGND VPWR VPWR _24730_/Q sky130_fd_sc_hd__dfrtp_4
X_21942_ _18314_/X VGND VGND VPWR VPWR _22027_/A sky130_fd_sc_hd__buf_2
XANTENNA__16589__B1 _16419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21873_ _16731_/Y VGND VGND VPWR VPWR _21879_/A sky130_fd_sc_hd__buf_2
X_24661_ _24169_/CLK _24661_/D HRESETn VGND VGND VPWR VPWR _24661_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_199_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23323__A1 _21881_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23323__B2 _21085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20698_/X _20823_/X _24927_/Q _20744_/A VGND VGND VPWR VPWR _24044_/D sky130_fd_sc_hd__a2bb2o_4
X_23612_ _23628_/CLK _23612_/D VGND VGND VPWR VPWR _23612_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24592_ _24592_/CLK _24592_/D HRESETn VGND VGND VPWR VPWR _15114_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20137__B2 _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20755_ _20739_/X _20754_/X _24911_/Q _20744_/X VGND VGND VPWR VPWR _20755_/X sky130_fd_sc_hd__a2bb2o_4
X_23543_ _23590_/CLK _20030_/X VGND VGND VPWR VPWR _23543_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12286__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23474_ _23514_/CLK _23474_/D VGND VGND VPWR VPWR _23474_/Q sky130_fd_sc_hd__dfxtp_4
X_20686_ _20686_/A _14291_/X VGND VGND VPWR VPWR _20686_/X sky130_fd_sc_hd__or2_4
XANTENNA__22429__A3 _22303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _15628_/Y _22425_/B VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__and2_4
X_25213_ _23385_/CLK _14213_/X HRESETn VGND VGND VPWR VPWR _20524_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22356_ _22352_/X _22355_/X _18306_/A VGND VGND VPWR VPWR _22356_/Y sky130_fd_sc_hd__o21ai_4
X_25144_ _25137_/CLK _25144_/D HRESETn VGND VGND VPWR VPWR _25144_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21307_ _24485_/Q _21307_/B VGND VGND VPWR VPWR _21307_/X sky130_fd_sc_hd__or2_4
X_25075_ _23690_/CLK _14718_/Y HRESETn VGND VGND VPWR VPWR _14683_/A sky130_fd_sc_hd__dfstp_4
X_22287_ _22283_/X _22285_/X _21308_/C _24831_/Q _22286_/X VGND VGND VPWR VPWR _22287_/X
+ sky130_fd_sc_hd__a32o_4
X_12040_ _25499_/Q VGND VGND VPWR VPWR _12040_/Y sky130_fd_sc_hd__inv_2
X_24026_ _24022_/CLK _20748_/X HRESETn VGND VGND VPWR VPWR _20746_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25549__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21238_ _21868_/B _21238_/B _21237_/X VGND VGND VPWR VPWR _21238_/X sky130_fd_sc_hd__and3_4
XFILLER_120_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21169_ _16548_/Y _21592_/A _21332_/A _21168_/X VGND VGND VPWR VPWR _21169_/X sky130_fd_sc_hd__a211o_4
XFILLER_238_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16221__A _24673_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23011__B1 _22816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13991_ _14028_/A VGND VGND VPWR VPWR _14027_/C sky130_fd_sc_hd__inv_2
XFILLER_105_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12302__B2 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15730_ _15726_/X VGND VGND VPWR VPWR _15730_/X sky130_fd_sc_hd__buf_2
X_12942_ _12944_/B VGND VGND VPWR VPWR _12942_/Y sky130_fd_sc_hd__inv_2
X_24928_ _24923_/CLK _24928_/D HRESETn VGND VGND VPWR VPWR _24928_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_207_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15661_ _21140_/A _17448_/C _15661_/C _13542_/C VGND VGND VPWR VPWR _15661_/X sky130_fd_sc_hd__or4_4
X_12873_ _12790_/Y _12878_/A _12872_/X VGND VGND VPWR VPWR _12873_/X sky130_fd_sc_hd__or3_4
X_24859_ _23386_/CLK _15785_/X HRESETn VGND VGND VPWR VPWR _21025_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18148__A _18051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17400_/A _17399_/X VGND VGND VPWR VPWR _17400_/X sky130_fd_sc_hd__or2_4
X_14612_ _14574_/B _14610_/Y _14608_/X _14611_/X _25093_/Q VGND VGND VPWR VPWR _25093_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11824_/A VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__inv_2
X_18380_ _18376_/Y _18379_/X _24202_/Q _18379_/X VGND VGND VPWR VPWR _18380_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15592_/A VGND VGND VPWR VPWR _15592_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A _17330_/X VGND VGND VPWR VPWR _17332_/C sky130_fd_sc_hd__nand2_4
XFILLER_199_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14543_ _14543_/A _14543_/B VGND VGND VPWR VPWR _14543_/X sky130_fd_sc_hd__and2_4
XANTENNA__20679__A2 _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ HWDATA[30] VGND VGND VPWR VPWR _11755_/X sky130_fd_sc_hd__buf_2
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17262_/A VGND VGND VPWR VPWR _17262_/Y sky130_fd_sc_hd__inv_2
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _14474_/A VGND VGND VPWR VPWR _14474_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11686_ _24236_/Q VGND VGND VPWR VPWR _11686_/Y sky130_fd_sc_hd__inv_2
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _19001_/A VGND VGND VPWR VPWR _19001_/Y sky130_fd_sc_hd__inv_2
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _16212_/Y _16210_/X _11773_/X _16210_/X VGND VGND VPWR VPWR _16213_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_197_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13425_ _13286_/X _23662_/Q VGND VGND VPWR VPWR _13425_/X sky130_fd_sc_hd__or2_4
X_17193_ _17193_/A VGND VGND VPWR VPWR _17193_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16143_/Y _16141_/X _11818_/X _16141_/X VGND VGND VPWR VPWR _16144_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13356_ _13356_/A _18949_/A VGND VGND VPWR VPWR _13358_/B sky130_fd_sc_hd__or2_4
XFILLER_6_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12307_ _25346_/Q _12305_/Y _13026_/C _24852_/Q VGND VGND VPWR VPWR _12307_/X sky130_fd_sc_hd__a2bb2o_4
X_16075_ _24725_/Q VGND VGND VPWR VPWR _16075_/Y sky130_fd_sc_hd__inv_2
X_13287_ _13286_/X _19681_/A VGND VGND VPWR VPWR _13287_/X sky130_fd_sc_hd__or2_4
XFILLER_216_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15026_ _15026_/A VGND VGND VPWR VPWR _15026_/Y sky130_fd_sc_hd__inv_2
X_19903_ _18282_/X _18285_/D _19481_/X VGND VGND VPWR VPWR _19904_/A sky130_fd_sc_hd__or3_4
X_12238_ _12503_/A VGND VGND VPWR VPWR _12238_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16807__B2 _16806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21800__A1 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ _25169_/Q _14347_/A _25167_/Q _12169_/D VGND VGND VPWR VPWR _12170_/B sky130_fd_sc_hd__and4_4
X_19834_ _23613_/Q VGND VGND VPWR VPWR _19834_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18272__A3 _15993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16977_ _17080_/A VGND VGND VPWR VPWR _17075_/C sky130_fd_sc_hd__inv_2
X_19765_ _19765_/A VGND VGND VPWR VPWR _19765_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14294__A1 _23444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19757__B1 _19734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20137__A2_N _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15970__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15928_ _15928_/A VGND VGND VPWR VPWR _15928_/Y sky130_fd_sc_hd__inv_2
X_18716_ _18715_/X VGND VGND VPWR VPWR _24161_/D sky130_fd_sc_hd__inv_2
X_19696_ _13162_/B VGND VGND VPWR VPWR _19696_/Y sky130_fd_sc_hd__inv_2
X_18647_ _24136_/Q VGND VGND VPWR VPWR _18648_/A sky130_fd_sc_hd__inv_2
X_15859_ _21045_/A _14462_/A VGND VGND VPWR VPWR _21173_/B sky130_fd_sc_hd__or2_4
XFILLER_91_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24854__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _18476_/A _18572_/B VGND VGND VPWR VPWR _18578_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17529_ _24298_/Q VGND VGND VPWR VPWR _17529_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20540_ _15465_/A _20540_/B _20682_/B VGND VGND VPWR VPWR _20540_/X sky130_fd_sc_hd__and3_4
XANTENNA__21212__A _21212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20471_ _20462_/X _20471_/B VGND VGND VPWR VPWR _20476_/B sky130_fd_sc_hd__and2_4
XANTENNA__16306__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22210_ _22210_/A _20153_/Y VGND VGND VPWR VPWR _22213_/B sky130_fd_sc_hd__or2_4
XFILLER_146_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23190_ _23148_/A VGND VGND VPWR VPWR _23190_/X sky130_fd_sc_hd__buf_2
XANTENNA__22292__A1 _22289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22292__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22141_ _15715_/X VGND VGND VPWR VPWR _22854_/B sky130_fd_sc_hd__buf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22072_ _22392_/A _22072_/B VGND VGND VPWR VPWR _22072_/X sky130_fd_sc_hd__or2_4
XFILLER_161_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23139__A _22479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23241__B1 _24291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21023_ _21023_/A _21023_/B VGND VGND VPWR VPWR _21023_/X sky130_fd_sc_hd__and2_4
XFILLER_102_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18263__A3 _15993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21882__A _21882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22974_ _12831_/Y _22725_/X _22861_/X _12593_/Y _22862_/X VGND VGND VPWR VPWR _22974_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__21555__B1 _25375_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24713_ _24697_/CLK _16109_/X HRESETn VGND VGND VPWR VPWR _23205_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17223__B2 _17322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21925_ _21895_/X _21925_/B VGND VGND VPWR VPWR _21925_/X sky130_fd_sc_hd__or2_4
XFILLER_16_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24595__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24644_ _24639_/CLK _24644_/D HRESETn VGND VGND VPWR VPWR _24644_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21856_ _16622_/A _21330_/X _21331_/X _21855_/X VGND VGND VPWR VPWR _21857_/C sky130_fd_sc_hd__a211o_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20788_/X _20806_/X _15583_/A _20792_/X VGND VGND VPWR VPWR _20807_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21787_ _21644_/A _21787_/B VGND VGND VPWR VPWR _21787_/X sky130_fd_sc_hd__or2_4
X_24575_ _24592_/CLK _24575_/D HRESETn VGND VGND VPWR VPWR _24575_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_125_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _25043_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19920__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23526_ _23597_/CLK _23526_/D VGND VGND VPWR VPWR _23526_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_188_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25215_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20738_ _20738_/A VGND VGND VPWR VPWR _20738_/Y sky130_fd_sc_hd__inv_2
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21122__A _21122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20669_ _17407_/B _20668_/Y _20669_/C VGND VGND VPWR VPWR _20669_/X sky130_fd_sc_hd__and3_4
X_23457_ _23454_/CLK _20266_/X VGND VGND VPWR VPWR _13313_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13182_/A VGND VGND VPWR VPWR _13315_/A sky130_fd_sc_hd__buf_2
X_22408_ _22408_/A _21656_/X VGND VGND VPWR VPWR _22408_/X sky130_fd_sc_hd__or2_4
X_14190_ _14190_/A _14131_/X VGND VGND VPWR VPWR _14190_/Y sky130_fd_sc_hd__nand2_4
X_23388_ _25365_/CLK HSEL VGND VGND VPWR VPWR _23351_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_152_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13141_ _13141_/A _13140_/X VGND VGND VPWR VPWR _13141_/X sky130_fd_sc_hd__or2_4
X_25127_ _25154_/CLK _14482_/X HRESETn VGND VGND VPWR VPWR _25127_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12771__B2 _24790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22339_ _22338_/Y _21353_/X _14227_/Y _14230_/A VGND VGND VPWR VPWR _22339_/X sky130_fd_sc_hd__o22a_4
XFILLER_152_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _12312_/X _13066_/B VGND VGND VPWR VPWR _13072_/Y sky130_fd_sc_hd__nand2_4
X_25058_ _23385_/CLK _14846_/X HRESETn VGND VGND VPWR VPWR _14826_/C sky130_fd_sc_hd__dfrtp_4
X_12023_ _25320_/Q VGND VGND VPWR VPWR _12023_/Y sky130_fd_sc_hd__inv_2
X_16900_ _16093_/Y _23332_/A _16093_/Y _23332_/A VGND VGND VPWR VPWR _16904_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24009_ _23980_/CLK _20688_/X HRESETn VGND VGND VPWR VPWR _24009_/Q sky130_fd_sc_hd__dfrtp_4
X_17880_ _16901_/Y _17877_/B VGND VGND VPWR VPWR _17880_/Y sky130_fd_sc_hd__nand2_4
XFILLER_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16831_ _14950_/Y _16828_/X HWDATA[17] _16828_/X VGND VGND VPWR VPWR _24436_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24216__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16598__A1_N _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15473__B1 _14420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19739__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19550_ _16464_/A _16464_/B _19550_/C _21382_/B VGND VGND VPWR VPWR _19551_/A sky130_fd_sc_hd__and4_4
X_16762_ _16762_/A VGND VGND VPWR VPWR _16762_/X sky130_fd_sc_hd__buf_2
XFILLER_219_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13974_ _14254_/A _13927_/X _14255_/A VGND VGND VPWR VPWR _13975_/B sky130_fd_sc_hd__or3_4
XFILLER_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18501_ _18488_/B _18499_/A VGND VGND VPWR VPWR _18502_/C sky130_fd_sc_hd__or2_4
X_15713_ _15751_/A VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__buf_2
X_12925_ _12819_/Y _12924_/X VGND VGND VPWR VPWR _12926_/B sky130_fd_sc_hd__or2_4
X_19481_ _17717_/X _24221_/Q _18288_/X VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__or3_4
XFILLER_74_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16693_ _16691_/Y _16692_/X _15752_/X _16692_/X VGND VGND VPWR VPWR _16693_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _16231_/A _18540_/B _16266_/Y _18434_/A VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15644_ _15643_/Y _15641_/X _15486_/X _15641_/X VGND VGND VPWR VPWR _15644_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_21_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12856_ _12783_/Y _12969_/A _12856_/C _12855_/X VGND VGND VPWR VPWR _12856_/X sky130_fd_sc_hd__or4_4
XPHY_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12638__B _12638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_84_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _25540_/Q VGND VGND VPWR VPWR _11807_/Y sky130_fd_sc_hd__inv_2
X_18363_ _18370_/A _18360_/Y _18362_/Y VGND VGND VPWR VPWR _18363_/X sky130_fd_sc_hd__a21o_4
XPHY_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15574_/Y _15572_/X _11758_/X _15572_/X VGND VGND VPWR VPWR _15575_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12787_ _25392_/Q VGND VGND VPWR VPWR _12787_/Y sky130_fd_sc_hd__inv_2
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17313_/X VGND VGND VPWR VPWR _24368_/D sky130_fd_sc_hd__inv_2
X_14526_ _14515_/Y VGND VGND VPWR VPWR _14526_/X sky130_fd_sc_hd__buf_2
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _24947_/Q _15515_/A _15517_/A _24944_/Q VGND VGND VPWR VPWR _11738_/X sky130_fd_sc_hd__or4_4
X_18294_ _18293_/X VGND VGND VPWR VPWR _18294_/X sky130_fd_sc_hd__buf_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13539__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23984__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17245_/A VGND VGND VPWR VPWR _17245_/Y sky130_fd_sc_hd__inv_2
X_14457_ _14446_/A VGND VGND VPWR VPWR _14457_/X sky130_fd_sc_hd__buf_2
X_11669_ _11668_/Y _22631_/A _11668_/Y _22631_/A VGND VGND VPWR VPWR _11675_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13209_/X _13392_/X _13407_/X _25334_/Q _13208_/A VGND VGND VPWR VPWR _13408_/X
+ sky130_fd_sc_hd__o32a_4
X_17176_ _16287_/Y _24377_/Q _16287_/Y _24377_/Q VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__a2bb2o_4
X_14388_ _14203_/X _14388_/B VGND VGND VPWR VPWR _14390_/B sky130_fd_sc_hd__or2_4
XFILLER_155_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16127_ _22920_/A VGND VGND VPWR VPWR _16127_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15965__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13339_ _13372_/A _23617_/Q VGND VGND VPWR VPWR _13340_/C sky130_fd_sc_hd__or2_4
XANTENNA__19437__A _19436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16058_ _24731_/Q VGND VGND VPWR VPWR _16058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15684__B _15683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15009_ _14973_/Y VGND VGND VPWR VPWR _15009_/X sky130_fd_sc_hd__buf_2
XANTENNA__13485__A _13484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17188__A2_N _17322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19817_ HWDATA[7] VGND VGND VPWR VPWR _19817_/X sky130_fd_sc_hd__buf_2
XANTENNA__18650__B1 _16601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16796__A _19131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19748_ _19742_/Y VGND VGND VPWR VPWR _19748_/X sky130_fd_sc_hd__buf_2
X_19679_ _19679_/A VGND VGND VPWR VPWR _19679_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21552__A3 _21550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21710_ _21530_/X _21709_/X _21445_/X _25528_/Q _22530_/B VGND VGND VPWR VPWR _21710_/X
+ sky130_fd_sc_hd__a32o_4
X_22690_ _20752_/Y _21123_/X _20891_/Y _21606_/X VGND VGND VPWR VPWR _22690_/X sky130_fd_sc_hd__o22a_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21641_ _21783_/A _20204_/Y VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__or2_4
XFILLER_197_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21572_ _21572_/A VGND VGND VPWR VPWR _21572_/Y sky130_fd_sc_hd__inv_2
X_24360_ _24346_/CLK _24360_/D HRESETn VGND VGND VPWR VPWR _24360_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12450__B1 _12403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20523_ _14286_/Y _20682_/B _24089_/Q VGND VGND VPWR VPWR _20527_/A sky130_fd_sc_hd__and3_4
X_23311_ _24550_/Q _22485_/X _22852_/X _23310_/X VGND VGND VPWR VPWR _23312_/C sky130_fd_sc_hd__a211o_4
XFILLER_166_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24291_ _24283_/CLK _17792_/Y HRESETn VGND VGND VPWR VPWR _24291_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20454_ _20613_/A _24095_/Q _20451_/X VGND VGND VPWR VPWR _20454_/X sky130_fd_sc_hd__o21a_4
X_23242_ _17243_/X _22493_/X _25401_/Q _22453_/X VGND VGND VPWR VPWR _23242_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23173_ _23208_/A _23161_/X _23173_/C _23172_/X VGND VGND VPWR VPWR _23173_/X sky130_fd_sc_hd__or4_4
XANTENNA__20815__A2 _20716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20385_ _20385_/A VGND VGND VPWR VPWR _20385_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22124_ _12238_/Y _15792_/X _16937_/Y _21457_/X VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22055_ _22055_/A _21976_/B VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__or2_4
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18236__A3 _18235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21776__B1 _14758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21006_ scl_oen_o_S5 _21005_/Y VGND VGND VPWR VPWR _21006_/X sky130_fd_sc_hd__and2_4
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24776__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23316__B _23313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24705__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22957_ _17229_/A _21065_/X VGND VGND VPWR VPWR _22960_/B sky130_fd_sc_hd__or2_4
XFILLER_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12710_ _12538_/Y _12710_/B VGND VGND VPWR VPWR _12737_/B sky130_fd_sc_hd__or2_4
X_21908_ _14700_/X VGND VGND VPWR VPWR _22373_/A sky130_fd_sc_hd__buf_2
XFILLER_216_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13690_ _13690_/A _13690_/B VGND VGND VPWR VPWR _13690_/X sky130_fd_sc_hd__or2_4
X_22888_ _17331_/A _22442_/A _12773_/A _22306_/X VGND VGND VPWR VPWR _22888_/X sky130_fd_sc_hd__a2bb2o_4
X_12641_ _12640_/X VGND VGND VPWR VPWR _25436_/D sky130_fd_sc_hd__inv_2
X_24627_ _24625_/CLK _16350_/X HRESETn VGND VGND VPWR VPWR _16348_/A sky130_fd_sc_hd__dfrtp_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23332__A _23332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21839_ _22400_/A _21839_/B _21839_/C VGND VGND VPWR VPWR _21839_/X sky130_fd_sc_hd__and3_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14954__A _14954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15360_ _15388_/A _15314_/X VGND VGND VPWR VPWR _15360_/X sky130_fd_sc_hd__or2_4
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12572_ _12572_/A VGND VGND VPWR VPWR _12572_/Y sky130_fd_sc_hd__inv_2
X_24558_ _24556_/CLK _16535_/X HRESETn VGND VGND VPWR VPWR _16532_/A sky130_fd_sc_hd__dfrtp_4
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16707__B1 _16609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21700__B1 _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _14308_/Y VGND VGND VPWR VPWR _14311_/X sky130_fd_sc_hd__buf_2
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23509_ _23493_/CLK _20125_/X VGND VGND VPWR VPWR _23509_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _15255_/X _15291_/B _15291_/C VGND VGND VPWR VPWR _15291_/X sky130_fd_sc_hd__and3_4
XFILLER_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24489_ _24493_/CLK _24489_/D HRESETn VGND VGND VPWR VPWR _24489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _17064_/A VGND VGND VPWR VPWR _17095_/A sky130_fd_sc_hd__buf_2
X_14242_ _25202_/Q VGND VGND VPWR VPWR _14242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21059__A2 _21039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14733__A2 _14713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14173_ _14153_/A _14172_/Y _25219_/Q _14153_/A VGND VGND VPWR VPWR _25219_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13124_ _13115_/X _13124_/B _13121_/C VGND VGND VPWR VPWR _25341_/D sky130_fd_sc_hd__and3_4
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18981_ _18981_/A VGND VGND VPWR VPWR _18981_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16903__A2_N _17752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12921__B _12819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22559__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11818__A _16245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13055_ _13055_/A VGND VGND VPWR VPWR _13055_/Y sky130_fd_sc_hd__inv_2
X_17932_ _24257_/Q _17931_/Y _17926_/X VGND VGND VPWR VPWR _17932_/X sky130_fd_sc_hd__o21a_4
X_12006_ _11999_/Y _12006_/B VGND VGND VPWR VPWR _12006_/Y sky130_fd_sc_hd__nor2_4
X_17863_ _24274_/Q _17863_/B VGND VGND VPWR VPWR _17865_/B sky130_fd_sc_hd__or2_4
XFILLER_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22411__A _22541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19602_ _19593_/Y _19601_/X _19439_/X _19601_/X VGND VGND VPWR VPWR _19602_/X sky130_fd_sc_hd__a2bb2o_4
X_16814_ _14914_/Y _16811_/X HWDATA[27] _16811_/X VGND VGND VPWR VPWR _16814_/X sky130_fd_sc_hd__a2bb2o_4
X_17794_ _17793_/X VGND VGND VPWR VPWR _17800_/B sky130_fd_sc_hd__inv_2
XFILLER_226_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15997__B2 _15947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16745_ _24479_/Q VGND VGND VPWR VPWR _16745_/Y sky130_fd_sc_hd__inv_2
X_19533_ _19533_/A VGND VGND VPWR VPWR _22039_/B sky130_fd_sc_hd__inv_2
XANTENNA__21027__A _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ _13943_/X VGND VGND VPWR VPWR _13957_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22731__A2 _22444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ _12908_/A _12908_/B _12907_/X VGND VGND VPWR VPWR _12908_/X sky130_fd_sc_hd__or3_4
X_19464_ _19463_/Y _19461_/X _19418_/X _19461_/X VGND VGND VPWR VPWR _23739_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19720__A _19719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16676_ _16675_/Y _16673_/X _16407_/X _16673_/X VGND VGND VPWR VPWR _24506_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13888_ _13880_/X _13887_/X _25192_/Q _13876_/A VGND VGND VPWR VPWR _25251_/D sky130_fd_sc_hd__o22a_4
XFILLER_34_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15627_ _15625_/Y _15621_/X _11838_/X _15626_/X VGND VGND VPWR VPWR _15627_/X sky130_fd_sc_hd__a2bb2o_4
X_18415_ _24660_/Q _18414_/A _16259_/Y _18476_/B VGND VGND VPWR VPWR _18415_/X sky130_fd_sc_hd__o22a_4
X_12839_ _25403_/Q VGND VGND VPWR VPWR _12839_/Y sky130_fd_sc_hd__inv_2
X_19395_ _19394_/Y _19392_/X _19305_/X _19392_/X VGND VGND VPWR VPWR _23763_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18346_ _18349_/B VGND VGND VPWR VPWR _18347_/B sky130_fd_sc_hd__inv_2
X_15558_ _11727_/A _15558_/B VGND VGND VPWR VPWR _15559_/D sky130_fd_sc_hd__or2_4
XFILLER_194_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14509_ _23970_/Q VGND VGND VPWR VPWR _14510_/C sky130_fd_sc_hd__inv_2
XFILLER_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18277_ _13789_/X VGND VGND VPWR VPWR _18277_/X sky130_fd_sc_hd__buf_2
XFILLER_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_171_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24101_/CLK sky130_fd_sc_hd__clkbuf_1
X_15489_ _16729_/A VGND VGND VPWR VPWR _15489_/X sky130_fd_sc_hd__buf_2
XFILLER_174_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17228_ _16363_/Y _17250_/A _24645_/Q _17227_/Y VGND VGND VPWR VPWR _17233_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_28_0_HCLK clkbuf_7_14_0_HCLK/X VGND VGND VPWR VPWR _25539_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17159_ _17159_/A _17159_/B VGND VGND VPWR VPWR _17160_/B sky130_fd_sc_hd__or2_4
XFILLER_128_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20170_ _19859_/X _13771_/X _18914_/X VGND VGND VPWR VPWR _20170_/X sky130_fd_sc_hd__or3_4
XFILLER_116_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12112__A1_N _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23860_ _23916_/CLK _23860_/D VGND VGND VPWR VPWR _13189_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22811_ _13607_/B _21967_/A _22706_/B _22527_/X VGND VGND VPWR VPWR _22811_/X sky130_fd_sc_hd__a211o_4
XFILLER_84_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12757__A1_N _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23791_ _23794_/CLK _19317_/X VGND VGND VPWR VPWR _13396_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22722__A2 _22425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25530_ _25528_/CLK _25530_/D HRESETn VGND VGND VPWR VPWR _25530_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22742_ _24434_/Q _22541_/X _22542_/X _22741_/X VGND VGND VPWR VPWR _22743_/C sky130_fd_sc_hd__a211o_4
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25461_ _25380_/CLK _25461_/D HRESETn VGND VGND VPWR VPWR _25461_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22673_ _22673_/A _22673_/B VGND VGND VPWR VPWR _22673_/X sky130_fd_sc_hd__or2_4
XFILLER_198_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24412_ _23926_/CLK _16895_/X HRESETn VGND VGND VPWR VPWR _20122_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21624_ _21617_/X _21623_/X _14721_/X VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22486__A1 _21881_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25392_ _25392_/CLK _12923_/X HRESETn VGND VGND VPWR VPWR _25392_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22486__B2 _22485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24343_ _24343_/CLK _24343_/D HRESETn VGND VGND VPWR VPWR _24343_/Q sky130_fd_sc_hd__dfstp_4
X_21555_ _17389_/A _21321_/X _25375_/Q _21535_/A VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22888__A1_N _17331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20506_ _23978_/Q _20683_/A VGND VGND VPWR VPWR _20506_/X sky130_fd_sc_hd__and2_4
X_21486_ _21482_/X _21485_/X _18306_/X VGND VGND VPWR VPWR _21487_/C sky130_fd_sc_hd__o21a_4
X_24274_ _24715_/CLK _17865_/X HRESETn VGND VGND VPWR VPWR _24274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20437_ _20437_/A _20437_/B VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__or2_4
X_23225_ _23188_/X _23222_/X _23224_/X VGND VGND VPWR VPWR _23226_/D sky130_fd_sc_hd__and3_4
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20368_ _20367_/Y _20365_/X _19629_/A _20365_/X VGND VGND VPWR VPWR _20368_/X sky130_fd_sc_hd__a2bb2o_4
X_23156_ _23156_/A _23146_/Y _23151_/X _23156_/D VGND VGND VPWR VPWR _23156_/X sky130_fd_sc_hd__or4_4
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22107_ _22107_/A _23274_/B VGND VGND VPWR VPWR _22111_/B sky130_fd_sc_hd__or2_4
X_23087_ _24576_/Q _23087_/B _22954_/C VGND VGND VPWR VPWR _23087_/X sky130_fd_sc_hd__and3_4
X_20299_ _23444_/Q _20298_/Y _23984_/Q _20297_/X VGND VGND VPWR VPWR _23444_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22038_ _21682_/A _22038_/B VGND VGND VPWR VPWR _22038_/X sky130_fd_sc_hd__or2_4
XFILLER_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22961__A2 _21456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ _14852_/X _14859_/Y _25054_/Q _14852_/X VGND VGND VPWR VPWR _14860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13811_ _25278_/Q VGND VGND VPWR VPWR _13811_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14791_ _14790_/X VGND VGND VPWR VPWR _14791_/X sky130_fd_sc_hd__buf_2
X_23989_ _24012_/CLK _20635_/Y HRESETn VGND VGND VPWR VPWR _17398_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22174__B1 _15676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16530_ _14420_/A VGND VGND VPWR VPWR _16530_/X sky130_fd_sc_hd__buf_2
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13742_ _13740_/B _13730_/X _13712_/X _13690_/B VGND VGND VPWR VPWR _25286_/D sky130_fd_sc_hd__o22a_4
XFILLER_217_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20686__A _20686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23062__A _22986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16461_ _22944_/A VGND VGND VPWR VPWR _22754_/A sky130_fd_sc_hd__buf_2
XFILLER_16_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13673_ _24070_/Q _20933_/B _13672_/X VGND VGND VPWR VPWR _13673_/X sky130_fd_sc_hd__or3_4
X_18200_ _18200_/A _23822_/Q VGND VGND VPWR VPWR _18200_/X sky130_fd_sc_hd__or2_4
XFILLER_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18156__A _13639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15600__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15412_ _15393_/A _15409_/B _15411_/Y VGND VGND VPWR VPWR _24989_/D sky130_fd_sc_hd__and3_4
X_12624_ _25407_/Q VGND VGND VPWR VPWR _12737_/A sky130_fd_sc_hd__inv_2
X_19180_ _19180_/A VGND VGND VPWR VPWR _19180_/Y sky130_fd_sc_hd__inv_2
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16392_ _15118_/Y _16384_/X _16389_/X _16391_/X VGND VGND VPWR VPWR _16392_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _18131_/A _18131_/B _18130_/X VGND VGND VPWR VPWR _18139_/B sky130_fd_sc_hd__or3_4
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15343_ _15357_/A _15343_/B _15342_/X VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__or3_4
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12555_ _24889_/Q VGND VGND VPWR VPWR _12555_/Y sky130_fd_sc_hd__inv_2
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_244_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _24989_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ _18165_/A _18062_/B VGND VGND VPWR VPWR _18063_/C sky130_fd_sc_hd__or2_4
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _15274_/A VGND VGND VPWR VPWR _15274_/Y sky130_fd_sc_hd__inv_2
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12229_/X _12212_/X _12480_/X VGND VGND VPWR VPWR _12486_/X sky130_fd_sc_hd__or3_4
XFILLER_8_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17013_ _16028_/Y _17018_/A _24731_/Q _17050_/D VGND VGND VPWR VPWR _17020_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14225_ _20686_/A VGND VGND VPWR VPWR _14225_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21310__A _15866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14156_ _14125_/A _14125_/B _14125_/A _14125_/B VGND VGND VPWR VPWR _14157_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18853__B1 _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13107_ _12386_/Y _13107_/B VGND VGND VPWR VPWR _13107_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24698__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14087_ _14066_/A VGND VGND VPWR VPWR _14087_/X sky130_fd_sc_hd__buf_2
X_18964_ _18963_/Y _18961_/X _17430_/X _18961_/X VGND VGND VPWR VPWR _23915_/D sky130_fd_sc_hd__a2bb2o_4
X_13038_ _13038_/A _13038_/B VGND VGND VPWR VPWR _13039_/B sky130_fd_sc_hd__or2_4
X_17915_ _17915_/A VGND VGND VPWR VPWR _17915_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18605__B1 _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24627__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _18876_/X _18890_/X _24127_/Q _24128_/Q _18893_/X VGND VGND VPWR VPWR _18895_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20412__B1 _11851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17846_ _17845_/X VGND VGND VPWR VPWR _24277_/D sky130_fd_sc_hd__inv_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20963__B2 _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14989_ _25019_/Q VGND VGND VPWR VPWR _15276_/A sky130_fd_sc_hd__inv_2
X_17777_ _23332_/A _17776_/Y VGND VGND VPWR VPWR _17779_/B sky130_fd_sc_hd__or2_4
XFILLER_207_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19516_ _21931_/B _19513_/X _11952_/X _19513_/X VGND VGND VPWR VPWR _23721_/D sky130_fd_sc_hd__a2bb2o_4
X_16728_ _24484_/Q VGND VGND VPWR VPWR _16728_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21912__B1 _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16659_ _16659_/A VGND VGND VPWR VPWR _23244_/A sky130_fd_sc_hd__inv_2
X_19447_ _19446_/Y _19444_/X _19377_/X _19444_/X VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_54_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _19376_/Y _19374_/X _19377_/X _19374_/X VGND VGND VPWR VPWR _23769_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18329_ _17464_/Y VGND VGND VPWR VPWR _20079_/A sky130_fd_sc_hd__buf_2
X_21340_ _21340_/A _22316_/B VGND VGND VPWR VPWR _21340_/X sky130_fd_sc_hd__or2_4
XANTENNA__14158__B1 _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22316__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21271_ _21271_/A _21271_/B VGND VGND VPWR VPWR _21272_/C sky130_fd_sc_hd__or2_4
XANTENNA__12842__A _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20222_ _21900_/B _20219_/X _19800_/A _20219_/X VGND VGND VPWR VPWR _23473_/D sky130_fd_sc_hd__a2bb2o_4
X_23010_ _24673_/Q _23010_/B VGND VGND VPWR VPWR _23013_/B sky130_fd_sc_hd__or2_4
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20153_ _20153_/A VGND VGND VPWR VPWR _20153_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19625__A _19624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20084_ _20083_/Y _20081_/X _19769_/X _20081_/X VGND VGND VPWR VPWR _23523_/D sky130_fd_sc_hd__a2bb2o_4
X_24961_ _23991_/CLK _15478_/X HRESETn VGND VGND VPWR VPWR _24961_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_112_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23912_ _24111_/CLK _23912_/D VGND VGND VPWR VPWR _13354_/B sky130_fd_sc_hd__dfxtp_4
X_24892_ _25062_/CLK _15708_/X HRESETn VGND VGND VPWR VPWR _24892_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20954__A1 _16662_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22986__A _22986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16083__B1 _15848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21890__A _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23843_ _23850_/CLK _19172_/X VGND VGND VPWR VPWR _23843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14919__D _14918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15830__B1 _24839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19021__B1 _18975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23774_ _23889_/CLK _19363_/X VGND VGND VPWR VPWR _18192_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _14408_/Y _14389_/X VGND VGND VPWR VPWR _23939_/D sky130_fd_sc_hd__and2_4
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25513_ _23555_/CLK _11945_/X HRESETn VGND VGND VPWR VPWR _19996_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22725_ _21316_/X VGND VGND VPWR VPWR _22725_/X sky130_fd_sc_hd__buf_2
XANTENNA__12439__D _12391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25444_ _25444_/CLK _12501_/X HRESETn VGND VGND VPWR VPWR _25444_/Q sky130_fd_sc_hd__dfrtp_4
X_22656_ _22655_/X VGND VGND VPWR VPWR _22656_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25206__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21607_ _21322_/A VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__buf_2
X_25375_ _24792_/CLK _25375_/D HRESETn VGND VGND VPWR VPWR _25375_/Q sky130_fd_sc_hd__dfrtp_4
X_22587_ _22586_/X VGND VGND VPWR VPWR _22587_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18704__A _18733_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12340_ _24834_/Q VGND VGND VPWR VPWR _12340_/Y sky130_fd_sc_hd__inv_2
X_24326_ _23534_/CLK _24326_/D HRESETn VGND VGND VPWR VPWR _24326_/Q sky130_fd_sc_hd__dfrtp_4
X_21538_ _21129_/X VGND VGND VPWR VPWR _21538_/X sky130_fd_sc_hd__buf_2
XFILLER_153_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12271_ _12262_/X _12265_/X _12267_/X _12270_/X VGND VGND VPWR VPWR _12281_/C sky130_fd_sc_hd__or4_4
X_24257_ _24258_/CLK _17932_/X HRESETn VGND VGND VPWR VPWR _24257_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19088__B1 _18991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_11_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23513_/CLK sky130_fd_sc_hd__clkbuf_1
X_21469_ _21468_/X _21469_/B VGND VGND VPWR VPWR _21469_/X sky130_fd_sc_hd__or2_4
XFILLER_181_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14010_ _25244_/Q _25243_/Q _14008_/X _14058_/C VGND VGND VPWR VPWR _14010_/X sky130_fd_sc_hd__or4_4
X_23208_ _23208_/A _23198_/X _23208_/C _23208_/D VGND VGND VPWR VPWR _23208_/X sky130_fd_sc_hd__or4_4
Xclkbuf_8_74_0_HCLK clkbuf_8_74_0_HCLK/A VGND VGND VPWR VPWR _24689_/CLK sky130_fd_sc_hd__clkbuf_1
X_24188_ _24194_/CLK _18519_/X HRESETn VGND VGND VPWR VPWR _24188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23139_ _22479_/A VGND VGND VPWR VPWR _23139_/X sky130_fd_sc_hd__buf_2
XFILLER_1_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24791__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15961_ _12268_/Y _15953_/X _15960_/X _15953_/X VGND VGND VPWR VPWR _24775_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24720__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14912_ _15074_/A VGND VGND VPWR VPWR _14912_/X sky130_fd_sc_hd__buf_2
X_17700_ _17701_/A _17701_/B VGND VGND VPWR VPWR _17700_/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15892_ _12774_/Y _15890_/X _11797_/X _15890_/X VGND VGND VPWR VPWR _24808_/D sky130_fd_sc_hd__a2bb2o_4
X_18680_ _18744_/A VGND VGND VPWR VPWR _18701_/A sky130_fd_sc_hd__inv_2
XFILLER_248_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16074__B1 _16073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14843_ _14826_/C _14811_/X _14826_/C _14811_/X VGND VGND VPWR VPWR _14843_/X sky130_fd_sc_hd__a2bb2o_4
X_17631_ _17591_/X _17610_/D _17553_/Y VGND VGND VPWR VPWR _17632_/C sky130_fd_sc_hd__o21a_4
XFILLER_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17562_ _17562_/A _17561_/X VGND VGND VPWR VPWR _17562_/X sky130_fd_sc_hd__or2_4
X_14774_ _13747_/A VGND VGND VPWR VPWR _14779_/A sky130_fd_sc_hd__buf_2
XANTENNA__22698__A1 _16284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11986_ _11981_/X _11985_/X VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__and2_4
X_16513_ _16533_/A VGND VGND VPWR VPWR _16513_/X sky130_fd_sc_hd__buf_2
X_19301_ _19301_/A VGND VGND VPWR VPWR _19301_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13725_ _13697_/A _13697_/B VGND VGND VPWR VPWR _13725_/Y sky130_fd_sc_hd__nand2_4
XFILLER_205_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17493_ _18335_/A _20079_/D VGND VGND VPWR VPWR _17494_/A sky130_fd_sc_hd__or2_4
XFILLER_210_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11831__A _11830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16444_ _15135_/Y _16442_/X _16073_/X _16442_/X VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__a2bb2o_4
X_19232_ _19232_/A VGND VGND VPWR VPWR _19232_/Y sky130_fd_sc_hd__inv_2
X_13656_ _25305_/Q _13649_/X _13655_/Y VGND VGND VPWR VPWR _13656_/X sky130_fd_sc_hd__o21a_4
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ _12607_/A _12602_/X _12603_/X _12607_/D VGND VGND VPWR VPWR _12608_/D sky130_fd_sc_hd__or4_4
X_19163_ _23845_/Q VGND VGND VPWR VPWR _19163_/Y sky130_fd_sc_hd__inv_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16729_/A VGND VGND VPWR VPWR _16375_/X sky130_fd_sc_hd__buf_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ _13587_/A _13580_/X _13587_/C _13586_/X VGND VGND VPWR VPWR _13587_/X sky130_fd_sc_hd__or4_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _17987_/A _18114_/B VGND VGND VPWR VPWR _18115_/C sky130_fd_sc_hd__or2_4
X_15326_ _15318_/X _15334_/D _15164_/Y VGND VGND VPWR VPWR _15327_/C sky130_fd_sc_hd__o21a_4
XFILLER_219_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12538_ _12538_/A VGND VGND VPWR VPWR _12538_/Y sky130_fd_sc_hd__inv_2
X_19094_ _19093_/Y _19090_/X _19048_/X _19090_/X VGND VGND VPWR VPWR _19094_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11858__A1_N _11853_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15888__B1 _11787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18045_ _17991_/X _18043_/X _18044_/X VGND VGND VPWR VPWR _18045_/X sky130_fd_sc_hd__and3_4
XANTENNA__21040__A _21032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15257_ _15071_/X _15256_/X VGND VGND VPWR VPWR _15257_/X sky130_fd_sc_hd__or2_4
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24879__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _12439_/B _12468_/X VGND VGND VPWR VPWR _12469_/X sky130_fd_sc_hd__or2_4
XANTENNA__12662__A _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14208_ _14207_/B _14205_/X _14209_/A VGND VGND VPWR VPWR _14208_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22622__A1 _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24808__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15188_ _15188_/A _15188_/B VGND VGND VPWR VPWR _15190_/B sky130_fd_sc_hd__or2_4
XFILLER_141_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14139_ _14141_/A _14136_/X _14137_/Y _14138_/X VGND VGND VPWR VPWR _14139_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19996_ _19996_/A VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__buf_2
XFILLER_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _23921_/Q VGND VGND VPWR VPWR _18947_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18878_ _23951_/Q _18877_/X VGND VGND VPWR VPWR _18878_/X sky130_fd_sc_hd__or2_4
XFILLER_228_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17829_ _16923_/Y _17834_/B _16964_/X VGND VGND VPWR VPWR _17829_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_243_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15812__B1 _11766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20840_ _16725_/Y _20833_/X _20836_/X _20839_/Y VGND VGND VPWR VPWR _20840_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21215__A _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20771_ _20776_/A VGND VGND VPWR VPWR _20772_/C sky130_fd_sc_hd__inv_2
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12837__A _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16309__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22510_ _22508_/X _22509_/X _22510_/C VGND VGND VPWR VPWR _22510_/X sky130_fd_sc_hd__or3_4
XANTENNA__11741__A _15661_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23490_ _24684_/CLK _23490_/D VGND VGND VPWR VPWR _23490_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_149_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23102__A2 _22851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18409__A1_N _24673_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22441_ _16354_/Y _22695_/B _22440_/X _16063_/Y _22283_/X VGND VGND VPWR VPWR _22442_/B
+ sky130_fd_sc_hd__o32a_4
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25160_ _25168_/CLK _14380_/X HRESETn VGND VGND VPWR VPWR _25160_/Q sky130_fd_sc_hd__dfrtp_4
X_22372_ _22095_/A _22372_/B VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__or2_4
X_24111_ _24111_/CLK MSI_S2 HRESETn VGND VGND VPWR VPWR _24111_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15879__B1 _11763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21323_ _17391_/A _21321_/X _13131_/A _21322_/X VGND VGND VPWR VPWR _21323_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20872__B1 _20863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25091_ _25276_/CLK _14616_/X HRESETn VGND VGND VPWR VPWR _13582_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12572__A _12572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21254_ _21271_/A _19116_/Y VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__or2_4
X_24042_ _24042_/CLK _20816_/Y HRESETn VGND VGND VPWR VPWR _24042_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24549__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20205_ _20193_/A VGND VGND VPWR VPWR _20205_/X sky130_fd_sc_hd__buf_2
X_21185_ _24217_/Q VGND VGND VPWR VPWR _21207_/A sky130_fd_sc_hd__buf_2
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20136_ _23505_/Q VGND VGND VPWR VPWR _21910_/B sky130_fd_sc_hd__inv_2
XFILLER_219_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _20067_/A VGND VGND VPWR VPWR _21922_/B sky130_fd_sc_hd__inv_2
X_24944_ _23408_/CLK _15521_/X HRESETn VGND VGND VPWR VPWR _24944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24875_ _24872_/CLK _15753_/X HRESETn VGND VGND VPWR VPWR _24875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15803__B1 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11840_ _25532_/Q VGND VGND VPWR VPWR _11840_/Y sky130_fd_sc_hd__inv_2
X_23826_ _23850_/CLK _23826_/D VGND VGND VPWR VPWR _18066_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11768_/Y _11769_/X _11770_/X _11769_/X VGND VGND VPWR VPWR _11771_/X sky130_fd_sc_hd__a2bb2o_4
X_23757_ _23735_/CLK _23757_/D VGND VGND VPWR VPWR _18207_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _25331_/Q _11712_/A _11979_/A VGND VGND VPWR VPWR _20969_/X sky130_fd_sc_hd__a21o_4
XANTENNA__17556__B1 _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13516_/A VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__buf_2
X_22708_ _22523_/X _22706_/X _21968_/A _22707_/Y VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__o22a_4
XFILLER_198_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14485_/A VGND VGND VPWR VPWR _14490_/X sky130_fd_sc_hd__buf_2
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _23703_/CLK _23688_/D VGND VGND VPWR VPWR _19610_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _13207_/A _13440_/X _25332_/Q _13267_/A VGND VGND VPWR VPWR _25332_/D sky130_fd_sc_hd__o22a_4
X_25427_ _25433_/CLK _12680_/X HRESETn VGND VGND VPWR VPWR _25427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23340__A _22810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22639_ _16601_/A _21067_/X _21755_/A _22638_/X VGND VGND VPWR VPWR _22639_/X sky130_fd_sc_hd__a211o_4
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16160_ _16159_/Y _16154_/X _16066_/X _16154_/X VGND VGND VPWR VPWR _24693_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13372_ _13372_/A _23616_/Q VGND VGND VPWR VPWR _13373_/C sky130_fd_sc_hd__or2_4
X_25358_ _25358_/CLK _13069_/X HRESETn VGND VGND VPWR VPWR _25358_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15111_ _24609_/Q VGND VGND VPWR VPWR _15111_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12323_ _25359_/Q VGND VGND VPWR VPWR _12323_/Y sky130_fd_sc_hd__inv_2
X_24309_ _24302_/CLK _24309_/D HRESETn VGND VGND VPWR VPWR _17666_/A sky130_fd_sc_hd__dfrtp_4
X_16091_ _11729_/X _15683_/X VGND VGND VPWR VPWR _16091_/X sky130_fd_sc_hd__or2_4
XANTENNA__24972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25289_ _24233_/CLK _25289_/D HRESETn VGND VGND VPWR VPWR _11678_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15042_ _15033_/X _15035_/X _15042_/C _15042_/D VGND VGND VPWR VPWR _15064_/A sky130_fd_sc_hd__or4_4
XFILLER_181_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14542__B1 _25119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12254_ _12424_/A _23049_/A _12424_/A _23049_/A VGND VGND VPWR VPWR _12260_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15885__A3 _15738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24901__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16889__A _14791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15793__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19850_ _19850_/A VGND VGND VPWR VPWR _19850_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _14338_/A _12182_/Y _11876_/X _12182_/Y VGND VGND VPWR VPWR _25470_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16295__B1 _16294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18801_ _18801_/A VGND VGND VPWR VPWR _24141_/D sky130_fd_sc_hd__inv_2
X_19781_ _19779_/Y _19780_/X _19734_/X _19780_/X VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16993_ _24730_/Q _24387_/Q _16060_/Y _16992_/Y VGND VGND VPWR VPWR _16993_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11826__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18732_ _18732_/A VGND VGND VPWR VPWR _18732_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15944_ _15938_/X _15943_/X HWDATA[30] _24783_/Q _15941_/X VGND VGND VPWR VPWR _24783_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16047__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15875_ _15896_/A VGND VGND VPWR VPWR _15875_/Y sky130_fd_sc_hd__inv_2
X_18663_ _24151_/Q VGND VGND VPWR VPWR _18696_/D sky130_fd_sc_hd__inv_2
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14826_ _14811_/C _14825_/X _14826_/C VGND VGND VPWR VPWR _14826_/X sky130_fd_sc_hd__or3_4
X_17614_ _17616_/B VGND VGND VPWR VPWR _17615_/B sky130_fd_sc_hd__inv_2
XFILLER_236_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18594_ _18595_/A _18598_/A VGND VGND VPWR VPWR _18594_/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21035__A _21035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14757_ _25068_/Q VGND VGND VPWR VPWR _22221_/A sky130_fd_sc_hd__buf_2
X_17545_ _11799_/Y _17535_/A _25546_/Q _17579_/A VGND VGND VPWR VPWR _17545_/X sky130_fd_sc_hd__a2bb2o_4
X_11969_ _11979_/B VGND VGND VPWR VPWR _11970_/D sky130_fd_sc_hd__inv_2
XANTENNA__12657__A _12657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _11705_/Y _13711_/B VGND VGND VPWR VPWR _13708_/X sky130_fd_sc_hd__or2_4
XFILLER_232_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17476_ _17478_/B VGND VGND VPWR VPWR _17477_/B sky130_fd_sc_hd__inv_2
XFILLER_220_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14688_ _21240_/A VGND VGND VPWR VPWR _14688_/X sky130_fd_sc_hd__buf_2
X_19215_ _19214_/Y _19212_/X _19148_/X _19212_/X VGND VGND VPWR VPWR _23827_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23250__A _23250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13639_ _25083_/Q VGND VGND VPWR VPWR _13639_/X sky130_fd_sc_hd__buf_2
X_16427_ _16427_/A VGND VGND VPWR VPWR _16427_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15968__A _15947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23096__B2 _21607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16358_ _24623_/Q VGND VGND VPWR VPWR _16358_/Y sky130_fd_sc_hd__inv_2
X_19146_ _19141_/Y _19145_/X _19032_/X _19145_/X VGND VGND VPWR VPWR _23852_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22843__B2 _22298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15309_ _24991_/Q VGND VGND VPWR VPWR _15407_/A sky130_fd_sc_hd__inv_2
XFILLER_145_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16289_ _16288_/X VGND VGND VPWR VPWR _16290_/A sky130_fd_sc_hd__buf_2
X_19077_ _19090_/A VGND VGND VPWR VPWR _19077_/X sky130_fd_sc_hd__buf_2
XANTENNA__12392__A _12391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18028_ _18069_/A _18028_/B _18027_/X VGND VGND VPWR VPWR _18028_/X sky130_fd_sc_hd__and3_4
XFILLER_160_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24642__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16799__A _24452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19979_ _19979_/A VGND VGND VPWR VPWR _19979_/X sky130_fd_sc_hd__buf_2
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22990_ _21129_/X VGND VGND VPWR VPWR _22990_/X sky130_fd_sc_hd__buf_2
XFILLER_228_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21941_ _21941_/A _20372_/Y VGND VGND VPWR VPWR _21945_/B sky130_fd_sc_hd__or2_4
XFILLER_216_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24660_ _24171_/CLK _24660_/D HRESETn VGND VGND VPWR VPWR _24660_/Q sky130_fd_sc_hd__dfrtp_4
X_21872_ _21872_/A _21868_/X _21871_/X VGND VGND VPWR VPWR _21872_/X sky130_fd_sc_hd__and3_4
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _25068_/CLK _23611_/D VGND VGND VPWR VPWR _23611_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_243_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20821_/Y _20818_/X _20822_/X VGND VGND VPWR VPWR _20823_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24591_ _24602_/CLK _24591_/D HRESETn VGND VGND VPWR VPWR _24591_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23542_ _23590_/CLK _20032_/X VGND VGND VPWR VPWR _20031_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_211_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20754_ _20752_/Y _20749_/Y _20753_/X VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__o21a_4
XFILLER_211_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _23577_/CLK _23473_/D VGND VGND VPWR VPWR _20221_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20685_ _20683_/A VGND VGND VPWR VPWR _20685_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_24_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25212_ _25212_/CLK _14215_/X HRESETn VGND VGND VPWR VPWR _14214_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21098__B1 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22424_ _16711_/Y _22424_/B VGND VGND VPWR VPWR _22424_/X sky130_fd_sc_hd__and2_4
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25143_ _25137_/CLK _25143_/D HRESETn VGND VGND VPWR VPWR _25143_/Q sky130_fd_sc_hd__dfstp_4
X_22355_ _21949_/A _22353_/X _22355_/C VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__and3_4
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21306_ _21306_/A VGND VGND VPWR VPWR _21320_/A sky130_fd_sc_hd__buf_2
XANTENNA__24383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25074_ _23690_/CLK _14733_/X HRESETn VGND VGND VPWR VPWR _13748_/A sky130_fd_sc_hd__dfrtp_4
X_22286_ _22425_/B VGND VGND VPWR VPWR _22286_/X sky130_fd_sc_hd__buf_2
XFILLER_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24025_ _24022_/CLK _20745_/X HRESETn VGND VGND VPWR VPWR _13139_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19085__A _19085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21237_ _21046_/X _21234_/X _21235_/X _21236_/Y VGND VGND VPWR VPWR _21237_/X sky130_fd_sc_hd__a211o_4
XFILLER_116_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16277__B1 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20073__B2 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21168_ _18515_/A _21173_/B _21173_/C VGND VGND VPWR VPWR _21168_/X sky130_fd_sc_hd__and3_4
XFILLER_172_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_148_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _25093_/CLK sky130_fd_sc_hd__clkbuf_1
X_20119_ _20119_/A VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__buf_2
XANTENNA__23011__A1 _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13990_ _14011_/A VGND VGND VPWR VPWR _14028_/A sky130_fd_sc_hd__buf_2
X_21099_ _23087_/B _21091_/X _21098_/X VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__and3_4
XFILLER_219_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16029__B1 _15960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ _12941_/A _12940_/X VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__or2_4
X_24927_ _24923_/CLK _15575_/X HRESETn VGND VGND VPWR VPWR _24927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_234_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13861__A _24007_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15660_ _15652_/Y _15655_/X _15656_/X _21026_/B _15659_/X VGND VGND VPWR VPWR _24897_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_206_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12872_ _12872_/A _12871_/X VGND VGND VPWR VPWR _12872_/X sky130_fd_sc_hd__or2_4
X_24858_ _23386_/CLK _24858_/D HRESETn VGND VGND VPWR VPWR _23386_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_34_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/A VGND VGND VPWR VPWR _14611_/X sky130_fd_sc_hd__buf_2
XANTENNA__23314__A2 _22673_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11820_/Y _11814_/X _11822_/X _11814_/X VGND VGND VPWR VPWR _25537_/D sky130_fd_sc_hd__a2bb2o_4
X_23809_ _23529_/CLK _23809_/D VGND VGND VPWR VPWR _23809_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15588_/Y _15584_/X _11780_/X _15590_/X VGND VGND VPWR VPWR _24921_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _25062_/CLK _24789_/D HRESETn VGND VGND VPWR VPWR _13548_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17330_/A _17330_/B VGND VGND VPWR VPWR _17330_/X sky130_fd_sc_hd__or2_4
XFILLER_14_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _23969_/Q _14541_/X _25119_/Q _14515_/Y VGND VGND VPWR VPWR _14542_/X sky130_fd_sc_hd__o22a_4
XPHY_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11754_/A VGND VGND VPWR VPWR _11754_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17341_/A _17338_/A _17322_/A _17229_/Y VGND VGND VPWR VPWR _17261_/X sky130_fd_sc_hd__or4_4
XFILLER_159_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23070__A _15588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14472_/Y _14468_/X _14412_/X _14468_/X VGND VGND VPWR VPWR _14473_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11685_/A VGND VGND VPWR VPWR _11685_/Y sky130_fd_sc_hd__inv_2
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16212_/A VGND VGND VPWR VPWR _16212_/Y sky130_fd_sc_hd__inv_2
X_19000_ _18998_/Y _14674_/A _18999_/X _14674_/A VGND VGND VPWR VPWR _23901_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ _13456_/A _13424_/B _13424_/C VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__and3_4
X_17192_ _24635_/Q _24364_/Q _16327_/Y _17331_/A VGND VGND VPWR VPWR _17200_/A sky130_fd_sc_hd__o22a_4
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16143_ _22673_/A VGND VGND VPWR VPWR _16143_/Y sky130_fd_sc_hd__inv_2
X_13355_ _13387_/A _13353_/X _13355_/C VGND VGND VPWR VPWR _13359_/B sky130_fd_sc_hd__and3_4
XFILLER_6_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _12306_/A VGND VGND VPWR VPWR _13026_/C sky130_fd_sc_hd__inv_2
XFILLER_155_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16074_ _16072_/Y _16069_/X _16073_/X _16069_/X VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__a2bb2o_4
X_13286_ _13228_/A VGND VGND VPWR VPWR _13286_/X sky130_fd_sc_hd__buf_2
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22414__A _23027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15025_ _15195_/A _15024_/Y _15292_/A _24452_/Q VGND VGND VPWR VPWR _15030_/B sky130_fd_sc_hd__a2bb2o_4
X_19902_ _23588_/Q VGND VGND VPWR VPWR _19902_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12237_ _24770_/Q VGND VGND VPWR VPWR _12237_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_44_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12940__A _12638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16412__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19833_ _19831_/Y _19829_/X _19832_/X _19829_/X VGND VGND VPWR VPWR _19833_/X sky130_fd_sc_hd__a2bb2o_4
X_12168_ _20982_/B VGND VGND VPWR VPWR _12168_/X sky130_fd_sc_hd__buf_2
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19206__B1 _19184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19764_ _18334_/X _18938_/B _18938_/C VGND VGND VPWR VPWR _19765_/A sky130_fd_sc_hd__or3_4
XANTENNA__16283__A3 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12099_ _12099_/A VGND VGND VPWR VPWR _12099_/Y sky130_fd_sc_hd__inv_2
X_16976_ _24399_/Q VGND VGND VPWR VPWR _17105_/A sky130_fd_sc_hd__inv_2
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14294__A2 _14289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18715_ _18678_/Y _18712_/X _18708_/B _18714_/X VGND VGND VPWR VPWR _18715_/X sky130_fd_sc_hd__a211o_4
XFILLER_110_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15927_ _15691_/X _15707_/X _15921_/X _15926_/X VGND VGND VPWR VPWR _15928_/A sky130_fd_sc_hd__a211o_4
X_19695_ _19694_/Y _19689_/X _19620_/X _19675_/Y VGND VGND VPWR VPWR _19695_/X sky130_fd_sc_hd__a2bb2o_4
X_18646_ _24132_/Q VGND VGND VPWR VPWR _18689_/C sky130_fd_sc_hd__inv_2
X_15858_ _15713_/X VGND VGND VPWR VPWR _15858_/X sky130_fd_sc_hd__buf_2
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16440__B1 _16157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14809_ _25052_/Q _14809_/B _14824_/A VGND VGND VPWR VPWR _14810_/B sky130_fd_sc_hd__or3_4
X_18577_ _18556_/X _18573_/X _18576_/Y VGND VGND VPWR VPWR _18577_/X sky130_fd_sc_hd__and3_4
X_15789_ _15561_/Y _15678_/X _15782_/X _13150_/A _15788_/X VGND VGND VPWR VPWR _24857_/D
+ sky130_fd_sc_hd__a32o_4
X_17528_ _25534_/Q _24305_/Q _11833_/Y _17684_/A VGND VGND VPWR VPWR _17533_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21867__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24894__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17459_ _17459_/A VGND VGND VPWR VPWR _18937_/B sky130_fd_sc_hd__buf_2
XANTENNA__24823__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20470_ _20470_/A _20470_/B VGND VGND VPWR VPWR _20471_/B sky130_fd_sc_hd__and2_4
XFILLER_118_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19129_ _19128_/Y _19126_/X _19085_/X _19126_/X VGND VGND VPWR VPWR _19129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22140_ _21547_/X _22139_/X _21550_/X _12572_/A _21551_/X VGND VGND VPWR VPWR _22140_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_146_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22071_ _22373_/A _22071_/B _22070_/X VGND VGND VPWR VPWR _22071_/X sky130_fd_sc_hd__and3_4
XANTENNA__19445__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23241__B2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21022_ _21071_/A _21022_/B VGND VGND VPWR VPWR _21022_/X sky130_fd_sc_hd__and2_4
XFILLER_141_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19633__A _19624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_1_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22973_ _23106_/A _22972_/X VGND VGND VPWR VPWR _22973_/Y sky130_fd_sc_hd__nor2_4
XFILLER_74_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21555__B2 _21535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24712_ _24712_/CLK _16112_/X HRESETn VGND VGND VPWR VPWR _24712_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21924_ _22093_/A _21924_/B VGND VGND VPWR VPWR _21926_/B sky130_fd_sc_hd__or2_4
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16431__B1 _16245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24643_ _24641_/CLK _24643_/D HRESETn VGND VGND VPWR VPWR _24643_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21855_ _24556_/Q _21855_/B _21752_/B VGND VGND VPWR VPWR _21855_/X sky130_fd_sc_hd__and3_4
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20804_/Y _20801_/Y _20809_/A VGND VGND VPWR VPWR _20806_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24574_ _24592_/CLK _24574_/D HRESETn VGND VGND VPWR VPWR _24574_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21786_ _21781_/X _21784_/X _21785_/X VGND VGND VPWR VPWR _21794_/B sky130_fd_sc_hd__o21a_4
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _23493_/CLK _20077_/X VGND VGND VPWR VPWR _20076_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20737_ _15623_/Y _20716_/X _20724_/X _20736_/X VGND VGND VPWR VPWR _20738_/A sky130_fd_sc_hd__o22a_4
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23454_/CLK _20268_/X VGND VGND VPWR VPWR _13350_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24564__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20668_ _20668_/A _17406_/B VGND VGND VPWR VPWR _20668_/Y sky130_fd_sc_hd__nand2_4
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22407_ _21996_/A _20344_/X VGND VGND VPWR VPWR _22407_/X sky130_fd_sc_hd__or2_4
XFILLER_137_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12220__A1 _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23387_ _24029_/CLK _20830_/A VGND VGND VPWR VPWR _23387_/Q sky130_fd_sc_hd__dfxtp_4
X_20599_ _20598_/X VGND VGND VPWR VPWR _20599_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16498__B1 _16412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _20746_/A _13139_/X VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__or2_4
X_25126_ _25125_/CLK _25126_/D HRESETn VGND VGND VPWR VPWR _25126_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20294__B2 _20291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22338_ _22338_/A VGND VGND VPWR VPWR _22338_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18855__A1_N _24569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13071_ _13069_/A _13068_/B _13071_/C VGND VGND VPWR VPWR _13071_/X sky130_fd_sc_hd__and3_4
X_25057_ _24343_/CLK _25057_/D HRESETn VGND VGND VPWR VPWR _14811_/C sky130_fd_sc_hd__dfrtp_4
X_22269_ _22265_/A _22267_/X _22268_/X VGND VGND VPWR VPWR _22269_/X sky130_fd_sc_hd__and3_4
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12022_ _11999_/Y _12006_/B _12006_/Y _12021_/X VGND VGND VPWR VPWR _12035_/A sky130_fd_sc_hd__a211o_4
X_24008_ _23976_/CLK _24008_/D HRESETn VGND VGND VPWR VPWR _24008_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16830_ _14922_/Y _16828_/X HWDATA[18] _16828_/X VGND VGND VPWR VPWR _24437_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16670__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19739__B2 _19719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13973_ _13940_/Y _14257_/D _13959_/X _15438_/C VGND VGND VPWR VPWR _14255_/A sky130_fd_sc_hd__or4_4
X_16761_ _24470_/Q VGND VGND VPWR VPWR _16761_/Y sky130_fd_sc_hd__inv_2
X_18500_ _24192_/Q _18500_/B VGND VGND VPWR VPWR _18500_/X sky130_fd_sc_hd__or2_4
XFILLER_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12924_ _12921_/C _12921_/D VGND VGND VPWR VPWR _12924_/X sky130_fd_sc_hd__or2_4
X_15712_ _15854_/B VGND VGND VPWR VPWR _15751_/A sky130_fd_sc_hd__inv_2
X_16692_ _16685_/A VGND VGND VPWR VPWR _16692_/X sky130_fd_sc_hd__buf_2
X_19480_ _20015_/B VGND VGND VPWR VPWR _19480_/X sky130_fd_sc_hd__buf_2
XFILLER_206_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18431_ _24180_/Q VGND VGND VPWR VPWR _18540_/B sky130_fd_sc_hd__inv_2
X_12855_ _12855_/A _12777_/A _12855_/C _12854_/X VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__or4_4
X_15643_ _15643_/A VGND VGND VPWR VPWR _15643_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17998__A _18006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15776__A2 _15774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11802_/Y _11804_/X _11805_/X _11804_/X VGND VGND VPWR VPWR _25541_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15574_ _24927_/Q VGND VGND VPWR VPWR _15574_/Y sky130_fd_sc_hd__inv_2
X_18362_ _18361_/X VGND VGND VPWR VPWR _18362_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12832__A2_N _23162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12786_ _12786_/A _12779_/X _12786_/C _12785_/X VGND VGND VPWR VPWR _12800_/C sky130_fd_sc_hd__or4_4
XPHY_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11798__B1 _11797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _20609_/A _14520_/X _25113_/Q _14522_/X VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__o22a_4
X_17313_ _17296_/A _17313_/B _17313_/C VGND VGND VPWR VPWR _17313_/X sky130_fd_sc_hd__or3_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21313__A _21300_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _24943_/Q _15524_/A VGND VGND VPWR VPWR _11737_/X sky130_fd_sc_hd__or2_4
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _18289_/C _17712_/A VGND VGND VPWR VPWR _18293_/X sky130_fd_sc_hd__or2_4
XANTENNA__16407__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13539__A1 _13526_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14455_/Y _14451_/X _14412_/X _14451_/X VGND VGND VPWR VPWR _25138_/D sky130_fd_sc_hd__a2bb2o_4
X_17244_ _17244_/A VGND VGND VPWR VPWR _17270_/C sky130_fd_sc_hd__inv_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _13702_/A VGND VGND VPWR VPWR _11668_/Y sky130_fd_sc_hd__inv_2
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13186_/Y _13399_/X _13406_/X VGND VGND VPWR VPWR _13407_/X sky130_fd_sc_hd__and3_4
X_17175_ _16345_/Y _24357_/Q _16345_/Y _24357_/Q VGND VGND VPWR VPWR _17181_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14387_ _14386_/X VGND VGND VPWR VPWR _14388_/B sky130_fd_sc_hd__buf_2
XFILLER_183_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16126_ _16125_/Y _16123_/X _15965_/X _16123_/X VGND VGND VPWR VPWR _24706_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16489__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13338_ _13371_/A _23633_/Q VGND VGND VPWR VPWR _13338_/X sky130_fd_sc_hd__or2_4
XFILLER_183_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20285__B2 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16690__A1_N _16689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18341__B _17459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ _16055_/Y _16056_/X _11827_/X _16056_/X VGND VGND VPWR VPWR _16057_/X sky130_fd_sc_hd__a2bb2o_4
X_13269_ _13211_/A VGND VGND VPWR VPWR _13412_/A sky130_fd_sc_hd__buf_2
XANTENNA__19427__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15008_ _14990_/X _24454_/Q _14990_/X _24454_/Q VGND VGND VPWR VPWR _15011_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20967__A1_N _20836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19816_ _19816_/A VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__buf_2
XFILLER_229_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_131_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23754_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16661__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19747_ _13297_/B VGND VGND VPWR VPWR _19747_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16959_ _16161_/Y _22199_/A _16169_/Y _24266_/Q VGND VGND VPWR VPWR _16959_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_194_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24169_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18069__A _18069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19678_ _19673_/Y _19676_/X _19677_/X _19676_/X VGND VGND VPWR VPWR _19678_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16413__B1 _16412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _16571_/A _24155_/Q _16571_/Y _18682_/A VGND VGND VPWR VPWR _18629_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21640_ _14766_/X VGND VGND VPWR VPWR _21783_/A sky130_fd_sc_hd__buf_2
XANTENNA__22319__A _22171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21571_ _14218_/Y _14202_/X _14244_/Y _14230_/A VGND VGND VPWR VPWR _21572_/A sky130_fd_sc_hd__o22a_4
XFILLER_177_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23310_ _16472_/A _23184_/X _23148_/X VGND VGND VPWR VPWR _23310_/X sky130_fd_sc_hd__o21a_4
X_20522_ _13982_/A _20519_/X _20521_/X VGND VGND VPWR VPWR _20522_/X sky130_fd_sc_hd__or3_4
XFILLER_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14727__B1 _14725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ _24272_/CLK _17797_/X HRESETn VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_177_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23241_ _12401_/B _21542_/X _24291_/Q _22501_/X VGND VGND VPWR VPWR _23241_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20453_ _24099_/Q _20451_/X VGND VGND VPWR VPWR _20455_/C sky130_fd_sc_hd__and2_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21877__B _21877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23172_ _23123_/X _23167_/Y _23168_/X _23171_/X VGND VGND VPWR VPWR _23172_/X sky130_fd_sc_hd__a2bb2o_4
X_20384_ _19527_/C _19986_/X _19505_/X VGND VGND VPWR VPWR _20385_/A sky130_fd_sc_hd__or3_4
XFILLER_173_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22123_ _22120_/X _22122_/X _21064_/X VGND VGND VPWR VPWR _22123_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22989__A _24638_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22054_ _22055_/A _21976_/B VGND VGND VPWR VPWR _22054_/X sky130_fd_sc_hd__and2_4
XFILLER_248_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21005_ _21005_/A VGND VGND VPWR VPWR _21005_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_90_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22956_ _23025_/A _22956_/B _22956_/C VGND VGND VPWR VPWR _22956_/X sky130_fd_sc_hd__and3_4
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16404__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21907_ _22380_/A _21907_/B _21907_/C VGND VGND VPWR VPWR _21907_/X sky130_fd_sc_hd__and3_4
XFILLER_244_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22887_ _12208_/Y _22507_/X _24281_/Q _21079_/A VGND VGND VPWR VPWR _22887_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16955__B2 _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12640_ _12633_/Y _12640_/B _12640_/C VGND VGND VPWR VPWR _12640_/X sky130_fd_sc_hd__or3_4
X_24626_ _24625_/CLK _16353_/X HRESETn VGND VGND VPWR VPWR _24626_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21838_ _13793_/D _21838_/B VGND VGND VPWR VPWR _21839_/C sky130_fd_sc_hd__or2_4
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24745__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _24861_/Q VGND VGND VPWR VPWR _12571_/Y sky130_fd_sc_hd__inv_2
X_24557_ _24556_/CLK _16538_/X HRESETn VGND VGND VPWR VPWR _24557_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21769_ _21765_/X _21768_/X _14721_/X VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__o21a_4
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12755__A _22302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17904__B1 _22003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _14310_/A _14305_/X _14310_/C VGND VGND VPWR VPWR _25185_/D sky130_fd_sc_hd__and3_4
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23508_ _24684_/CLK _20130_/X VGND VGND VPWR VPWR _20126_/A sky130_fd_sc_hd__dfxtp_4
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18172__A3 _18171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15131__A _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15290_ _15290_/A _15293_/B VGND VGND VPWR VPWR _15291_/C sky130_fd_sc_hd__nand2_4
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24488_ _24488_/CLK _24488_/D HRESETn VGND VGND VPWR VPWR _24488_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _14240_/Y _14238_/X _13806_/X _14238_/X VGND VGND VPWR VPWR _14241_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23439_ _23553_/CLK _23439_/D VGND VGND VPWR VPWR _23439_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14172_ _14138_/X _14171_/X _25139_/Q _14141_/A VGND VGND VPWR VPWR _14172_/Y sky130_fd_sc_hd__a22oi_4
X_13123_ _13003_/A _13123_/B VGND VGND VPWR VPWR _13124_/B sky130_fd_sc_hd__or2_4
X_25109_ _23970_/CLK _25109_/D HRESETn VGND VGND VPWR VPWR _21560_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_180_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18980_ _18979_/Y _18974_/X _17452_/X _18974_/A VGND VGND VPWR VPWR _18980_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _13054_/A _13053_/X VGND VGND VPWR VPWR _13055_/A sky130_fd_sc_hd__or2_4
X_17931_ _17930_/X VGND VGND VPWR VPWR _17931_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12005_ _24107_/Q _12002_/X _12004_/Y VGND VGND VPWR VPWR _12006_/B sky130_fd_sc_hd__o21a_4
X_17862_ _17864_/B VGND VGND VPWR VPWR _17863_/B sky130_fd_sc_hd__inv_2
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19601_ _19615_/A VGND VGND VPWR VPWR _19601_/X sky130_fd_sc_hd__buf_2
X_16813_ _14976_/Y _16811_/X HWDATA[28] _16811_/X VGND VGND VPWR VPWR _16813_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21308__A _21320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17793_ _17609_/B _17793_/B VGND VGND VPWR VPWR _17793_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_204_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24552_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_219_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23226__C _23221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19532_ _22245_/B _19529_/X _11943_/X _19529_/X VGND VGND VPWR VPWR _23715_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11834__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16744_ _15014_/Y _16739_/X _16389_/X _16743_/X VGND VGND VPWR VPWR _24480_/D sky130_fd_sc_hd__a2bb2o_4
X_13956_ _15435_/B _13955_/X VGND VGND VPWR VPWR _13956_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14210__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17199__A1 _24624_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17199__B2 _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12907_ _12895_/B _12871_/X _12825_/Y VGND VGND VPWR VPWR _12907_/X sky130_fd_sc_hd__o21a_4
X_19463_ _19463_/A VGND VGND VPWR VPWR _19463_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13887_ _21568_/A _13869_/X _25250_/Q _13864_/X VGND VGND VPWR VPWR _13887_/X sky130_fd_sc_hd__o22a_4
X_16675_ _24506_/Q VGND VGND VPWR VPWR _16675_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12771__A2_N _24790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18414_ _18414_/A VGND VGND VPWR VPWR _18476_/B sky130_fd_sc_hd__inv_2
XFILLER_50_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12838_ _12837_/Y _21712_/A _12853_/A _12804_/Y VGND VGND VPWR VPWR _12838_/X sky130_fd_sc_hd__a2bb2o_4
X_15626_ _15626_/A VGND VGND VPWR VPWR _15626_/X sky130_fd_sc_hd__buf_2
XANTENNA__24486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19394_ _19394_/A VGND VGND VPWR VPWR _19394_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22139__A _22139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18345_ _11661_/A _18333_/B _17485_/Y VGND VGND VPWR VPWR _18349_/B sky130_fd_sc_hd__o21a_4
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _12857_/A _12767_/Y _12888_/A _12768_/Y VGND VGND VPWR VPWR _12772_/C sky130_fd_sc_hd__a2bb2o_4
X_15557_ _15758_/A VGND VGND VPWR VPWR _15557_/X sky130_fd_sc_hd__buf_2
XANTENNA__19896__B1 _19643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _23395_/Q _20461_/C _14506_/X _25118_/Q _14507_/Y VGND VGND VPWR VPWR _14508_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _14885_/Y _15485_/X _14479_/X _15485_/X VGND VGND VPWR VPWR _24957_/D sky130_fd_sc_hd__a2bb2o_4
X_18276_ _13804_/D _18262_/X _13481_/A _23360_/A _18269_/X VGND VGND VPWR VPWR _24226_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_187_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15083__A2_N _16434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17227_ _24374_/Q VGND VGND VPWR VPWR _17227_/Y sky130_fd_sc_hd__inv_2
X_14439_ _25143_/Q VGND VGND VPWR VPWR _14439_/Y sky130_fd_sc_hd__inv_2
X_17158_ _17139_/B VGND VGND VPWR VPWR _17159_/B sky130_fd_sc_hd__inv_2
XFILLER_155_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16109_ _16108_/Y _16104_/X _15952_/X _16104_/X VGND VGND VPWR VPWR _16109_/X sky130_fd_sc_hd__a2bb2o_4
X_17089_ _17037_/Y _17088_/X _17065_/X VGND VGND VPWR VPWR _17089_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21758__A1 _21606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__19820__B1 _19769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22810_ _22810_/A _22809_/X VGND VGND VPWR VPWR _22810_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__11744__A _21332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23790_ _23794_/CLK _19319_/X VGND VGND VPWR VPWR _13428_/B sky130_fd_sc_hd__dfxtp_4
X_22741_ _16770_/A _22543_/X _22544_/X VGND VGND VPWR VPWR _22741_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_240_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25460_ _25380_/CLK _12437_/Y HRESETn VGND VGND VPWR VPWR _25460_/Q sky130_fd_sc_hd__dfrtp_4
X_22672_ _22155_/B VGND VGND VPWR VPWR _22673_/B sky130_fd_sc_hd__buf_2
XFILLER_241_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24411_ _25068_/CLK _16898_/X HRESETn VGND VGND VPWR VPWR _20146_/A sky130_fd_sc_hd__dfrtp_4
X_21623_ _21646_/A _21623_/B _21622_/X VGND VGND VPWR VPWR _21623_/X sky130_fd_sc_hd__and3_4
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25391_ _25392_/CLK _25391_/D HRESETn VGND VGND VPWR VPWR _12773_/A sky130_fd_sc_hd__dfrtp_4
X_24342_ _24343_/CLK _17417_/X HRESETn VGND VGND VPWR VPWR _21008_/A sky130_fd_sc_hd__dfstp_4
XFILLER_194_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21554_ _12232_/Y _21542_/A _16929_/A _21440_/X VGND VGND VPWR VPWR _21554_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20505_ _20493_/X _20505_/B VGND VGND VPWR VPWR _20505_/X sky130_fd_sc_hd__or2_4
X_24273_ _24272_/CLK _24273_/D HRESETn VGND VGND VPWR VPWR _24273_/Q sky130_fd_sc_hd__dfrtp_4
X_21485_ _21485_/A _21483_/X _21484_/X VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__and3_4
XFILLER_165_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23224_ _14914_/A _22153_/X _23015_/X _23223_/X VGND VGND VPWR VPWR _23224_/X sky130_fd_sc_hd__a211o_4
X_20436_ _15495_/X VGND VGND VPWR VPWR _20437_/B sky130_fd_sc_hd__inv_2
X_23155_ _22950_/A _23152_/X _23154_/X VGND VGND VPWR VPWR _23156_/D sky130_fd_sc_hd__and3_4
X_20367_ _23418_/Q VGND VGND VPWR VPWR _20367_/Y sky130_fd_sc_hd__inv_2
X_22106_ _23009_/A VGND VGND VPWR VPWR _23253_/A sky130_fd_sc_hd__buf_2
XFILLER_121_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23086_ _16214_/A _22827_/B VGND VGND VPWR VPWR _23089_/B sky130_fd_sc_hd__or2_4
X_20298_ _20297_/X VGND VGND VPWR VPWR _20298_/Y sky130_fd_sc_hd__inv_2
X_22037_ _22033_/X _22036_/X _21697_/X VGND VGND VPWR VPWR _22037_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13810_ _13808_/Y _13805_/X _13809_/X _13805_/X VGND VGND VPWR VPWR _13810_/X sky130_fd_sc_hd__a2bb2o_4
X_14790_ _14789_/Y _14790_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__and2_4
XANTENNA__24926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23988_ _24012_/CLK _23988_/D HRESETn VGND VGND VPWR VPWR _20627_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_180_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22174__A1 _16617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13741_ _13690_/X _13740_/X _13689_/X _13722_/X _11691_/A VGND VGND VPWR VPWR _25287_/D
+ sky130_fd_sc_hd__a32o_4
X_22939_ _16226_/A _23010_/B VGND VGND VPWR VPWR _22939_/X sky130_fd_sc_hd__or2_4
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16928__A1 _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_34_0_HCLK clkbuf_8_34_0_HCLK/A VGND VGND VPWR VPWR _23628_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_204_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_18_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ _13672_/A _13671_/X _24062_/Q _24061_/Q VGND VGND VPWR VPWR _13672_/X sky130_fd_sc_hd__or4_4
X_16460_ _16460_/A VGND VGND VPWR VPWR _22944_/A sky130_fd_sc_hd__buf_2
XFILLER_188_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_97_0_HCLK clkbuf_8_97_0_HCLK/A VGND VGND VPWR VPWR _24642_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12623_ _12740_/A _12742_/A _12623_/C _12623_/D VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__or4_4
X_15411_ _15411_/A _15401_/X VGND VGND VPWR VPWR _15411_/Y sky130_fd_sc_hd__nand2_4
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16391_ _16415_/A VGND VGND VPWR VPWR _16391_/X sky130_fd_sc_hd__buf_2
X_24609_ _24602_/CLK _16404_/X HRESETn VGND VGND VPWR VPWR _24609_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15342_ _15316_/X _15334_/D _15096_/Y VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__o21a_4
X_18130_ _18130_/A _18128_/X _18130_/C VGND VGND VPWR VPWR _18130_/X sky130_fd_sc_hd__and3_4
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12554_ _12644_/A VGND VGND VPWR VPWR _12631_/C sky130_fd_sc_hd__inv_2
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20075__A2_N _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _15268_/A _15259_/X _14996_/X _15270_/B VGND VGND VPWR VPWR _15274_/A sky130_fd_sc_hd__a211o_4
X_18061_ _18008_/A VGND VGND VPWR VPWR _18165_/A sky130_fd_sc_hd__buf_2
X_12485_ _12501_/A _12485_/B _12485_/C VGND VGND VPWR VPWR _25449_/D sky130_fd_sc_hd__and3_4
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__B1 SCLK_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14224_ _21004_/A _14219_/X _13819_/X _14210_/A VGND VGND VPWR VPWR _25208_/D sky130_fd_sc_hd__a2bb2o_4
X_17012_ _17008_/X _17012_/B _17010_/X _17011_/X VGND VGND VPWR VPWR _17026_/B sky130_fd_sc_hd__or4_4
X_14155_ _14141_/A VGND VGND VPWR VPWR _14155_/X sky130_fd_sc_hd__buf_2
XANTENNA__11829__A _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13106_ _13104_/A _13106_/B _13105_/Y VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__and3_4
X_14086_ _14013_/B _14074_/X _14066_/X _14013_/A _14085_/X VGND VGND VPWR VPWR _25242_/D
+ sky130_fd_sc_hd__a32o_4
X_18963_ _18963_/A VGND VGND VPWR VPWR _18963_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13037_ _12992_/Y _13052_/B _12370_/Y _12999_/X VGND VGND VPWR VPWR _13038_/B sky130_fd_sc_hd__or4_4
X_17914_ _17907_/A _17907_/B VGND VGND VPWR VPWR _17914_/X sky130_fd_sc_hd__or2_4
X_18894_ _18876_/X _18890_/X _24128_/Q _24129_/Q _18893_/X VGND VGND VPWR VPWR _24129_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16616__B1 _16530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21038__A _22947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17845_ _17766_/B _17818_/X _17790_/X _17842_/B VGND VGND VPWR VPWR _17845_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24667__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ _17776_/A VGND VGND VPWR VPWR _17776_/Y sky130_fd_sc_hd__inv_2
X_14988_ _15002_/A _14976_/Y _15258_/A _24423_/Q VGND VGND VPWR VPWR _14988_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19515_ _23721_/Q VGND VGND VPWR VPWR _21931_/B sky130_fd_sc_hd__inv_2
X_16727_ _16725_/Y _16721_/X _16726_/X _16721_/X VGND VGND VPWR VPWR _24485_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13939_ _13931_/Y _13932_/X _13935_/X _13948_/C VGND VGND VPWR VPWR _13940_/A sky130_fd_sc_hd__or4_4
XFILLER_208_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16919__B2 _17753_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13850__B1 _13849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17251__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19446_ _18081_/B VGND VGND VPWR VPWR _19446_/Y sky130_fd_sc_hd__inv_2
X_16658_ _16657_/Y _16655_/X _16389_/X _16655_/X VGND VGND VPWR VPWR _24513_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15609_ _15614_/A VGND VGND VPWR VPWR _15609_/X sky130_fd_sc_hd__buf_2
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_5_0_HCLK clkbuf_5_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19377_ _19085_/A VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__buf_2
X_16589_ _16588_/Y _16584_/X _16419_/X _16584_/X VGND VGND VPWR VPWR _16589_/X sky130_fd_sc_hd__a2bb2o_4
X_18328_ _21834_/A _18327_/Y _17901_/Y VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18541__B1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18259_ _11670_/Y _18258_/X _17430_/X _18258_/X VGND VGND VPWR VPWR _24237_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22316__B _22316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21270_ _21273_/A _20295_/Y VGND VGND VPWR VPWR _21272_/B sky130_fd_sc_hd__or2_4
XFILLER_156_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20221_ _20221_/A VGND VGND VPWR VPWR _21900_/B sky130_fd_sc_hd__inv_2
XFILLER_143_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16855__B1 _16537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20152_ _20148_/Y _20151_/X _20102_/X _20151_/X VGND VGND VPWR VPWR _20152_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22928__B1 _25392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24960_ _23991_/CLK _15481_/X HRESETn VGND VGND VPWR VPWR _15479_/A sky130_fd_sc_hd__dfstp_4
X_20083_ _23523_/Q VGND VGND VPWR VPWR _20083_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16607__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20403__B2 _20385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23911_ _24111_/CLK _23911_/D VGND VGND VPWR VPWR _18973_/A sky130_fd_sc_hd__dfxtp_4
X_24891_ _24825_/CLK _15721_/X HRESETn VGND VGND VPWR VPWR _24891_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20954__A2 _20854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23842_ _23830_/CLK _19175_/X VGND VGND VPWR VPWR _18062_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23773_ _23850_/CLK _19365_/X VGND VGND VPWR VPWR _18224_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19276__A2_N _19271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_250_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _24340_/CLK sky130_fd_sc_hd__clkbuf_1
X_20985_ _20463_/A _22115_/A _14550_/A VGND VGND VPWR VPWR _23936_/D sky130_fd_sc_hd__a21o_4
XANTENNA__13841__B1 _11834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22724_ _22724_/A _21868_/B VGND VGND VPWR VPWR _22724_/X sky130_fd_sc_hd__or2_4
X_25512_ _23441_/CLK _11949_/X HRESETn VGND VGND VPWR VPWR _20000_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_225_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23105__B1 _12330_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25443_ _25443_/CLK _25443_/D HRESETn VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22655_ _21063_/A _22650_/X _21844_/X _22654_/Y VGND VGND VPWR VPWR _22655_/X sky130_fd_sc_hd__a211o_4
XFILLER_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21606_ _21606_/A VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__buf_2
X_25374_ _24799_/CLK _25374_/D HRESETn VGND VGND VPWR VPWR _12853_/A sky130_fd_sc_hd__dfrtp_4
X_22586_ _22567_/Y _22573_/Y _22582_/Y _21455_/X _22585_/X VGND VGND VPWR VPWR _22586_/X
+ sky130_fd_sc_hd__a32o_4
X_24325_ _24327_/CLK _17608_/X HRESETn VGND VGND VPWR VPWR _17525_/A sky130_fd_sc_hd__dfrtp_4
X_21537_ _21537_/A _21536_/X VGND VGND VPWR VPWR _21537_/X sky130_fd_sc_hd__or2_4
XANTENNA__23972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12270_ _25460_/Q _12268_/Y _12269_/Y _24773_/Q VGND VGND VPWR VPWR _12270_/X sky130_fd_sc_hd__a2bb2o_4
X_24256_ _24258_/CLK _24256_/D HRESETn VGND VGND VPWR VPWR _13550_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_153_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21130__B _21046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21468_ _22271_/A VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__buf_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15543__A2_N _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23207_ _23123_/X _23204_/Y _23168_/X _23206_/X VGND VGND VPWR VPWR _23208_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20419_ _20996_/B _20419_/B VGND VGND VPWR VPWR _20419_/X sky130_fd_sc_hd__or2_4
X_24187_ _23973_/CLK _18521_/X HRESETn VGND VGND VPWR VPWR _24187_/Q sky130_fd_sc_hd__dfrtp_4
X_21399_ _21398_/X _19295_/Y VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__or2_4
XFILLER_108_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23138_ _16666_/Y _23177_/B VGND VGND VPWR VPWR _23138_/X sky130_fd_sc_hd__and2_4
XANTENNA__23338__A _22535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20106__A1_N _20104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24341__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15960_ HWDATA[22] VGND VGND VPWR VPWR _15960_/X sky130_fd_sc_hd__buf_2
X_23069_ _16671_/Y _23177_/B VGND VGND VPWR VPWR _23069_/X sky130_fd_sc_hd__and2_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14679__B _14679_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14911_ _25023_/Q _14909_/Y _14910_/Y _24445_/Q VGND VGND VPWR VPWR _14911_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15891_ _12788_/Y _15887_/X _11793_/X _15890_/X VGND VGND VPWR VPWR _24809_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_60_0_HCLK clkbuf_5_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17630_ _17598_/A _17626_/B _17630_/C VGND VGND VPWR VPWR _17630_/X sky130_fd_sc_hd__and3_4
X_14842_ _24005_/D _14841_/X _20672_/A _24005_/D VGND VGND VPWR VPWR _25059_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24760__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17561_ _17542_/X _17561_/B _17555_/X _17561_/D VGND VGND VPWR VPWR _17561_/X sky130_fd_sc_hd__or4_4
XFILLER_63_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _11985_/A _11984_/X VGND VGND VPWR VPWR _11985_/X sky130_fd_sc_hd__and2_4
X_14773_ _14772_/X VGND VGND VPWR VPWR _14773_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13832__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19300_ _18937_/B _18905_/D _18334_/X _20256_/D VGND VGND VPWR VPWR _19301_/A sky130_fd_sc_hd__or4_4
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16512_ _16512_/A VGND VGND VPWR VPWR _16512_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13724_ _13699_/B _13716_/X _13721_/Y _13723_/X _11700_/A VGND VGND VPWR VPWR _25295_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17492_ _17486_/X VGND VGND VPWR VPWR _17492_/X sky130_fd_sc_hd__buf_2
X_19231_ _19230_/Y _19225_/X _19139_/X _19225_/A VGND VGND VPWR VPWR _23821_/D sky130_fd_sc_hd__a2bb2o_4
X_16443_ _15086_/Y _16442_/X _16070_/X _16442_/X VGND VGND VPWR VPWR _24591_/D sky130_fd_sc_hd__a2bb2o_4
X_13655_ _25305_/Q _14320_/A _13654_/X VGND VGND VPWR VPWR _13655_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__15585__B1 _11773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12729_/A _24866_/Q _12740_/A _24863_/Q VGND VGND VPWR VPWR _12607_/D sky130_fd_sc_hd__a2bb2o_4
X_19162_ _19161_/Y _19159_/X _19048_/X _19159_/X VGND VGND VPWR VPWR _19162_/X sky130_fd_sc_hd__a2bb2o_4
X_13586_ _25268_/Q _25096_/Q _13584_/Y _14603_/A VGND VGND VPWR VPWR _13586_/X sky130_fd_sc_hd__o22a_4
X_16374_ _24617_/Q VGND VGND VPWR VPWR _16374_/Y sky130_fd_sc_hd__inv_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ _18039_/A _23784_/Q VGND VGND VPWR VPWR _18115_/B sky130_fd_sc_hd__or2_4
X_12537_ _25427_/Q _12535_/Y _25433_/Q _12536_/Y VGND VGND VPWR VPWR _12537_/X sky130_fd_sc_hd__a2bb2o_4
X_15325_ _15337_/A _15294_/A VGND VGND VPWR VPWR _15334_/D sky130_fd_sc_hd__and2_4
X_19093_ _23870_/Q VGND VGND VPWR VPWR _19093_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18044_ _18178_/A _18044_/B VGND VGND VPWR VPWR _18044_/X sky130_fd_sc_hd__or2_4
X_12468_ _12292_/X _13017_/B VGND VGND VPWR VPWR _12468_/X sky130_fd_sc_hd__or2_4
X_15256_ _15256_/A _15172_/X VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__or2_4
X_14207_ _14816_/A _14207_/B VGND VGND VPWR VPWR _14209_/A sky130_fd_sc_hd__nor2_4
X_15187_ _15186_/X VGND VGND VPWR VPWR _15188_/B sky130_fd_sc_hd__inv_2
X_12399_ _12391_/X _12282_/X VGND VGND VPWR VPWR _12400_/B sky130_fd_sc_hd__and2_4
XANTENNA__22622__A2 _22678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16837__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14138_ _14132_/B VGND VGND VPWR VPWR _14138_/X sky130_fd_sc_hd__buf_2
XFILLER_140_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19995_ _23554_/Q VGND VGND VPWR VPWR _22047_/B sky130_fd_sc_hd__inv_2
XFILLER_140_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14069_ _14069_/A _14069_/B VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__or2_4
X_18946_ _18944_/Y _18940_/X _17433_/X _18945_/X VGND VGND VPWR VPWR _23922_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16150__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24848__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18877_ _20552_/A _20555_/B VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__or2_4
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24126__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17828_ _16914_/Y _17832_/A _17768_/D _17820_/B VGND VGND VPWR VPWR _17834_/B sky130_fd_sc_hd__or4_4
XANTENNA__19461__A _19460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _17758_/Y _16929_/Y _17759_/C VGND VGND VPWR VPWR _17759_/X sky130_fd_sc_hd__or3_4
XFILLER_63_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20770_ _20761_/X _20769_/X _24914_/Q _20765_/X VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__a2bb2o_4
X_19429_ _19415_/A VGND VGND VPWR VPWR _19429_/X sky130_fd_sc_hd__buf_2
XFILLER_223_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_80_0_HCLK clkbuf_7_40_0_HCLK/X VGND VGND VPWR VPWR _25402_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22440_ _22543_/A VGND VGND VPWR VPWR _22440_/X sky130_fd_sc_hd__buf_2
XFILLER_149_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ _22392_/A _22371_/B VGND VGND VPWR VPWR _22371_/X sky130_fd_sc_hd__or2_4
XFILLER_175_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24110_ _25316_/CLK _12035_/C HRESETn VGND VGND VPWR VPWR _12029_/A sky130_fd_sc_hd__dfrtp_4
X_21322_ _21322_/A VGND VGND VPWR VPWR _21322_/X sky130_fd_sc_hd__buf_2
XFILLER_164_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_HCLK clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR clkbuf_3_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_25090_ _25276_/CLK _25090_/D HRESETn VGND VGND VPWR VPWR _13575_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24041_ _24042_/CLK _20812_/X HRESETn VGND VGND VPWR VPWR _13127_/B sky130_fd_sc_hd__dfrtp_4
X_21253_ _21257_/A _21253_/B VGND VGND VPWR VPWR _21253_/X sky130_fd_sc_hd__or2_4
XANTENNA__19636__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20204_ _20204_/A VGND VGND VPWR VPWR _20204_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23158__A _24779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21184_ _17714_/A VGND VGND VPWR VPWR _21204_/A sky130_fd_sc_hd__inv_2
XFILLER_116_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20135_ _20133_/Y _20129_/X _20108_/X _20134_/X VGND VGND VPWR VPWR _23506_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17156__A _17064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24589__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20066_ _22086_/B _20060_/X _19796_/X _20065_/X VGND VGND VPWR VPWR _20066_/X sky130_fd_sc_hd__a2bb2o_4
X_24943_ _23408_/CLK _15523_/X HRESETn VGND VGND VPWR VPWR _24943_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24874_ _24872_/CLK _15755_/X HRESETn VGND VGND VPWR VPWR _24874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_234_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23825_ _23830_/CLK _19221_/X VGND VGND VPWR VPWR _18104_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_233_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13814__B1 _13812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ HWDATA[26] VGND VGND VPWR VPWR _11770_/X sky130_fd_sc_hd__buf_2
X_23756_ _25082_/CLK _19416_/X VGND VGND VPWR VPWR _19412_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_214_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20830_/A _13677_/A _13676_/X _24515_/Q _20883_/A VGND VGND VPWR VPWR _24078_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _22707_/A _22468_/X VGND VGND VPWR VPWR _22707_/Y sky130_fd_sc_hd__nor2_4
XFILLER_241_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23687_ _23703_/CLK _23687_/D VGND VGND VPWR VPWR _19614_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ _20878_/X _20898_/X _24498_/Q _20883_/X VGND VGND VPWR VPWR _20899_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13209_/A _13424_/X _13439_/X _25333_/Q _13208_/A VGND VGND VPWR VPWR _13440_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__25377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22638_ _16517_/A _22440_/X _22545_/X VGND VGND VPWR VPWR _22638_/X sky130_fd_sc_hd__o21a_4
X_25426_ _25433_/CLK _25426_/D HRESETn VGND VGND VPWR VPWR _25426_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_108_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24913_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13371_ _13371_/A _13371_/B VGND VGND VPWR VPWR _13373_/B sky130_fd_sc_hd__or2_4
X_25357_ _25358_/CLK _13071_/X HRESETn VGND VGND VPWR VPWR _25357_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13859__A _24008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22569_ _21129_/X VGND VGND VPWR VPWR _22569_/X sky130_fd_sc_hd__buf_2
XFILLER_186_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12322_ _12322_/A _12316_/X _12322_/C _12321_/X VGND VGND VPWR VPWR _12349_/B sky130_fd_sc_hd__or4_4
X_15110_ _25005_/Q VGND VGND VPWR VPWR _15347_/A sky130_fd_sc_hd__inv_2
XFILLER_6_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16090_ _13818_/A VGND VGND VPWR VPWR _16090_/X sky130_fd_sc_hd__buf_2
X_24308_ _24302_/CLK _24308_/D HRESETn VGND VGND VPWR VPWR _17581_/A sky130_fd_sc_hd__dfrtp_4
X_25288_ _24233_/CLK _13739_/X HRESETn VGND VGND VPWR VPWR _11702_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15041_ _25030_/Q _15039_/Y _15260_/C _15032_/A VGND VGND VPWR VPWR _15042_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12253_ _25461_/Q VGND VGND VPWR VPWR _12424_/A sky130_fd_sc_hd__inv_2
X_24239_ _24240_/CLK _24239_/D HRESETn VGND VGND VPWR VPWR _24239_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16819__B1 _15734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20615__A1 _20609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23068__A _23066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12184_ _12184_/A VGND VGND VPWR VPWR _14338_/A sky130_fd_sc_hd__inv_2
XANTENNA__15793__B _15792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18800_ _18794_/C _18799_/X _18729_/X _18795_/Y VGND VGND VPWR VPWR _18801_/A sky130_fd_sc_hd__a211o_4
X_19780_ _19765_/Y VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__buf_2
XANTENNA__24941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16992_ _24387_/Q VGND VGND VPWR VPWR _16992_/Y sky130_fd_sc_hd__inv_2
X_18731_ _18729_/X _18725_/Y _18731_/C VGND VGND VPWR VPWR _18732_/A sky130_fd_sc_hd__or3_4
X_15943_ _15863_/X VGND VGND VPWR VPWR _15943_/X sky130_fd_sc_hd__buf_2
XFILLER_77_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18662_ _16622_/Y _24135_/Q _16562_/A _18670_/A VGND VGND VPWR VPWR _18662_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15874_ _15858_/X _15865_/X _15723_/X _23290_/A _15872_/X VGND VGND VPWR VPWR _24820_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_225_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17613_ _17613_/A VGND VGND VPWR VPWR _17613_/Y sky130_fd_sc_hd__inv_2
X_14825_ _25055_/Q _14824_/X _25056_/Q VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__or3_4
X_18593_ _18425_/Y _18597_/B VGND VGND VPWR VPWR _18598_/A sky130_fd_sc_hd__or2_4
XFILLER_236_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16809__A2_N _16806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17544_ _11779_/Y _24319_/Q _11779_/Y _24319_/Q VGND VGND VPWR VPWR _17544_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14756_ _14725_/X _14755_/X _14725_/X _14755_/X VGND VGND VPWR VPWR _14756_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21035__B _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11968_ _11979_/A _11979_/B VGND VGND VPWR VPWR _11968_/X sky130_fd_sc_hd__or2_4
X_13707_ _11668_/Y _13707_/B VGND VGND VPWR VPWR _13711_/B sky130_fd_sc_hd__or2_4
X_17475_ _24213_/Q VGND VGND VPWR VPWR _17477_/A sky130_fd_sc_hd__inv_2
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11899_ _11883_/Y _11898_/B _25524_/Q _11898_/Y VGND VGND VPWR VPWR _25524_/D sky130_fd_sc_hd__o22a_4
X_14687_ _14687_/A VGND VGND VPWR VPWR _21275_/A sky130_fd_sc_hd__buf_2
XFILLER_205_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_67_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19214_ _19214_/A VGND VGND VPWR VPWR _19214_/Y sky130_fd_sc_hd__inv_2
X_16426_ _16425_/Y _16423_/X _16238_/X _16423_/X VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13638_ _25083_/Q VGND VGND VPWR VPWR _18089_/A sky130_fd_sc_hd__inv_2
XANTENNA__23096__A2 _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22147__A _22986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _19159_/A VGND VGND VPWR VPWR _19145_/X sky130_fd_sc_hd__buf_2
X_16357_ _16356_/Y _16352_/X _16066_/X _16352_/X VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__a2bb2o_4
X_13569_ _25099_/Q VGND VGND VPWR VPWR _14581_/A sky130_fd_sc_hd__inv_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12673__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23967__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15308_ _15120_/Y _15411_/A _15401_/A _15415_/A VGND VGND VPWR VPWR _15308_/X sky130_fd_sc_hd__or4_4
XFILLER_146_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19076_ _19075_/X VGND VGND VPWR VPWR _19090_/A sky130_fd_sc_hd__inv_2
X_16288_ _22513_/B _16288_/B VGND VGND VPWR VPWR _16288_/X sky130_fd_sc_hd__and2_4
X_18027_ _18027_/A _18027_/B _18026_/X VGND VGND VPWR VPWR _18027_/X sky130_fd_sc_hd__or3_4
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15239_ _15238_/X VGND VGND VPWR VPWR _25029_/D sky130_fd_sc_hd__inv_2
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16286__A1 _15678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19978_ _19978_/A VGND VGND VPWR VPWR _21675_/B sky130_fd_sc_hd__inv_2
XFILLER_141_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24682__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18929_ _18916_/Y VGND VGND VPWR VPWR _18929_/X sky130_fd_sc_hd__buf_2
XANTENNA__24611__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
X_21940_ _21934_/X _21939_/X _17732_/A VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__o21a_4
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21871_ _24725_/Q _22424_/B _21121_/A _21870_/X VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__a211o_4
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23610_ _23628_/CLK _23610_/D VGND VGND VPWR VPWR _19843_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11752__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20822_ _20822_/A _20822_/B _13145_/X VGND VGND VPWR VPWR _20822_/X sky130_fd_sc_hd__or3_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24590_ _24602_/CLK _16444_/X HRESETn VGND VGND VPWR VPWR _15135_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _23565_/CLK _20035_/X VGND VGND VPWR VPWR _20033_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_211_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16949__A1_N _16166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ _20752_/A _13141_/X VGND VGND VPWR VPWR _20753_/X sky130_fd_sc_hd__or2_4
XFILLER_223_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _23529_/CLK _20224_/X VGND VGND VPWR VPWR _20223_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ _20684_/A VGND VGND VPWR VPWR _20684_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25211_ _25212_/CLK _14217_/X HRESETn VGND VGND VPWR VPWR _20497_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22423_ _22294_/A _22422_/Y VGND VGND VPWR VPWR _22435_/C sky130_fd_sc_hd__nor2_4
XFILLER_137_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19160__B1 _19091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25142_ _25148_/CLK _14447_/X HRESETn VGND VGND VPWR VPWR _25142_/Q sky130_fd_sc_hd__dfstp_4
X_22354_ _21948_/A _22354_/B VGND VGND VPWR VPWR _22355_/C sky130_fd_sc_hd__or2_4
XFILLER_136_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21305_ _15650_/X VGND VGND VPWR VPWR _21306_/A sky130_fd_sc_hd__inv_2
XFILLER_124_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25073_ _25062_/CLK _14746_/X HRESETn VGND VGND VPWR VPWR _25073_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15894__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22285_ _22285_/A _22284_/X VGND VGND VPWR VPWR _22285_/X sky130_fd_sc_hd__or2_4
XFILLER_105_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22598__A1 _17362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24024_ _24495_/CLK _20738_/Y HRESETn VGND VGND VPWR VPWR _24024_/Q sky130_fd_sc_hd__dfrtp_4
X_21236_ _25304_/Q _21046_/X VGND VGND VPWR VPWR _21236_/Y sky130_fd_sc_hd__nor2_4
XFILLER_105_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21167_ _21167_/A _21172_/B VGND VGND VPWR VPWR _21170_/B sky130_fd_sc_hd__or2_4
X_20118_ _20100_/Y VGND VGND VPWR VPWR _20118_/X sky130_fd_sc_hd__buf_2
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21098_ _21047_/X _21095_/X _21096_/X _21097_/X VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__a211o_4
XFILLER_218_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17226__B1 _16348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12940_ _12638_/B _12856_/X VGND VGND VPWR VPWR _12940_/X sky130_fd_sc_hd__or2_4
X_20049_ _21807_/B _20044_/X _20003_/X _20044_/X VGND VGND VPWR VPWR _23536_/D sky130_fd_sc_hd__a2bb2o_4
X_24926_ _24923_/CLK _15578_/X HRESETn VGND VGND VPWR VPWR _24926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23335__B _16552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21136__A _21161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12871_ _12609_/X _12846_/X VGND VGND VPWR VPWR _12871_/X sky130_fd_sc_hd__and2_4
X_24857_ _23386_/CLK _24857_/D HRESETn VGND VGND VPWR VPWR _13150_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12758__A _12899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/A _14610_/B VGND VGND VPWR VPWR _14610_/Y sky130_fd_sc_hd__nand2_4
XFILLER_215_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11822_ _16248_/A VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__buf_2
X_23808_ _23529_/CLK _23808_/D VGND VGND VPWR VPWR _23808_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25558__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15614_/A VGND VGND VPWR VPWR _15590_/X sky130_fd_sc_hd__buf_2
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _24258_/CLK _15930_/X HRESETn VGND VGND VPWR VPWR _15920_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__21325__A2 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__B _12391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11715_/Y _11751_/X _11752_/X _11751_/X VGND VGND VPWR VPWR _25556_/D sky130_fd_sc_hd__a2bb2o_4
X_14541_ _25107_/Q _14519_/X _23395_/Q _14514_/X VGND VGND VPWR VPWR _14541_/X sky130_fd_sc_hd__o22a_4
XFILLER_199_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23739_ _23794_/CLK _23739_/D VGND VGND VPWR VPWR _19463_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_242_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _24360_/Q VGND VGND VPWR VPWR _17338_/A sky130_fd_sc_hd__inv_2
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11677_/X _11684_/B _11684_/C _11684_/D VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__or4_4
X_14472_ _25130_/Q VGND VGND VPWR VPWR _14472_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15788__B _15683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16209_/Y _16210_/X _11770_/X _16210_/X VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _13423_/A _13423_/B _13423_/C VGND VGND VPWR VPWR _13424_/C sky130_fd_sc_hd__or3_4
X_25409_ _25410_/CLK _25409_/D HRESETn VGND VGND VPWR VPWR _12599_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14763__A1 _21630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17191_ _24364_/Q VGND VGND VPWR VPWR _17331_/A sky130_fd_sc_hd__inv_2
XFILLER_127_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13354_ _13450_/A _13354_/B VGND VGND VPWR VPWR _13355_/C sky130_fd_sc_hd__or2_4
X_16142_ _16140_/Y _16136_/X _11813_/X _16141_/X VGND VGND VPWR VPWR _24700_/D sky130_fd_sc_hd__a2bb2o_4
X_12305_ _24831_/Q VGND VGND VPWR VPWR _12305_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13285_ _13285_/A _13285_/B _13285_/C VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__and3_4
X_16073_ _14427_/A VGND VGND VPWR VPWR _16073_/X sky130_fd_sc_hd__buf_2
XANTENNA__18180__A _18051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14722__A1_N _14721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12236_ _12236_/A _12207_/X _12236_/C _12235_/X VGND VGND VPWR VPWR _12282_/A sky130_fd_sc_hd__or4_4
X_15024_ _24478_/Q VGND VGND VPWR VPWR _15024_/Y sky130_fd_sc_hd__inv_2
X_19901_ _19899_/Y _19895_/X _19900_/X _19895_/A VGND VGND VPWR VPWR _23589_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_9_0_HCLK clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19832_ HWDATA[1] VGND VGND VPWR VPWR _19832_/X sky130_fd_sc_hd__buf_2
X_12167_ _14342_/B VGND VGND VPWR VPWR _20982_/B sky130_fd_sc_hd__buf_2
X_19763_ _13179_/B VGND VGND VPWR VPWR _19763_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12097_/Y _12095_/X _11871_/X _12095_/X VGND VGND VPWR VPWR _12098_/X sky130_fd_sc_hd__a2bb2o_4
X_16975_ _24731_/Q _17050_/D _16018_/Y _24404_/Q VGND VGND VPWR VPWR _16980_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18714_ _18714_/A VGND VGND VPWR VPWR _18714_/X sky130_fd_sc_hd__buf_2
XANTENNA__17217__B1 _24622_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15926_ _13597_/X _15703_/A _15923_/X _15925_/Y VGND VGND VPWR VPWR _15926_/X sky130_fd_sc_hd__a211o_4
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19694_ _13457_/B VGND VGND VPWR VPWR _19694_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22761__A1 _21307_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_30_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18645_ _24537_/Q _18764_/A _16620_/Y _24136_/Q VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__a2bb2o_4
X_15857_ _15678_/X _15713_/X _15851_/X _12989_/A _15856_/X VGND VGND VPWR VPWR _15857_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15779__B1 _15486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14808_ _14822_/C _14822_/B _14823_/A VGND VGND VPWR VPWR _14809_/B sky130_fd_sc_hd__or3_4
XANTENNA__25299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18576_ _18479_/D _18573_/B VGND VGND VPWR VPWR _18576_/Y sky130_fd_sc_hd__nand2_4
X_15788_ _15560_/X _15683_/X VGND VGND VPWR VPWR _15788_/X sky130_fd_sc_hd__or2_4
X_17527_ _24305_/Q VGND VGND VPWR VPWR _17684_/A sky130_fd_sc_hd__inv_2
XANTENNA__25228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14739_ _14736_/Y _14717_/X _14738_/Y VGND VGND VPWR VPWR _14739_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_177_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17458_ _24328_/Q _17455_/X _17458_/C VGND VGND VPWR VPWR _17459_/A sky130_fd_sc_hd__or3_4
XFILLER_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16409_ _16415_/A VGND VGND VPWR VPWR _16409_/X sky130_fd_sc_hd__buf_2
X_17389_ _17389_/A _17389_/B VGND VGND VPWR VPWR _17389_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15951__B1 _15950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19128_ _23857_/Q VGND VGND VPWR VPWR _19128_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20827__A1 _20825_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_154_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _23615_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22292__A3 _21308_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22605__A _22605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14506__A1 _14550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19059_ _19058_/Y _19056_/X _19008_/X _19056_/X VGND VGND VPWR VPWR _23883_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24863__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22070_ _22094_/A _22070_/B VGND VGND VPWR VPWR _22070_/X sky130_fd_sc_hd__or2_4
XFILLER_142_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21021_ _21021_/A _21109_/A VGND VGND VPWR VPWR _23378_/A sky130_fd_sc_hd__and2_4
XFILLER_248_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22972_ _12266_/Y _22286_/X _22730_/X _12375_/Y _22858_/X VGND VGND VPWR VPWR _22972_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__23155__B _23152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24711_ _24712_/CLK _16114_/X HRESETn VGND VGND VPWR VPWR _24711_/Q sky130_fd_sc_hd__dfrtp_4
X_21923_ _22235_/A _21923_/B _21922_/X VGND VGND VPWR VPWR _21923_/X sky130_fd_sc_hd__and3_4
X_21854_ _16268_/A _22945_/A VGND VGND VPWR VPWR _21857_/B sky130_fd_sc_hd__or2_4
X_24642_ _24642_/CLK _24642_/D HRESETn VGND VGND VPWR VPWR _16308_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15785__A3 _15782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22504__B2 _16003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20805_ _13145_/A _13145_/B _13144_/X VGND VGND VPWR VPWR _20809_/A sky130_fd_sc_hd__or3_4
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21251_/X VGND VGND VPWR VPWR _21785_/X sky130_fd_sc_hd__buf_2
X_24573_ _24537_/CLK _16496_/X HRESETn VGND VGND VPWR VPWR _24573_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20735_/Y _20731_/X _13138_/X VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__o21a_4
X_23524_ _23522_/CLK _23524_/D VGND VGND VPWR VPWR _23524_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_50_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23454_/CLK _23455_/D VGND VGND VPWR VPWR _23455_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20667_ _20667_/A VGND VGND VPWR VPWR _20667_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22406_ _22406_/A VGND VGND VPWR VPWR _22406_/Y sky130_fd_sc_hd__inv_2
X_23386_ _23386_/CLK _23386_/D VGND VGND VPWR VPWR _23386_/Q sky130_fd_sc_hd__dfxtp_4
X_20598_ _14430_/Y _20550_/Y _20564_/X _20597_/X VGND VGND VPWR VPWR _20598_/X sky130_fd_sc_hd__a211o_4
XFILLER_192_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22337_ _14816_/A _21733_/B _20681_/A _22190_/B VGND VGND VPWR VPWR _22337_/X sky130_fd_sc_hd__a2bb2o_4
X_25125_ _25125_/CLK _25125_/D HRESETn VGND VGND VPWR VPWR _14487_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_192_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ _13063_/B _13066_/X VGND VGND VPWR VPWR _13071_/C sky130_fd_sc_hd__nand2_4
X_25056_ _24343_/CLK _14853_/X HRESETn VGND VGND VPWR VPWR _25056_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22268_ _22264_/A _22268_/B VGND VGND VPWR VPWR _22268_/X sky130_fd_sc_hd__or2_4
XANTENNA__24533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12021_ _12011_/X _12012_/X _12021_/C _12020_/X VGND VGND VPWR VPWR _12021_/X sky130_fd_sc_hd__or4_4
X_24007_ _23976_/CLK _24007_/D HRESETn VGND VGND VPWR VPWR _24007_/Q sky130_fd_sc_hd__dfrtp_4
X_21219_ _18268_/A _21216_/X _21218_/X _23360_/A _13802_/A VGND VGND VPWR VPWR _21220_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_104_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22199_ _22199_/A _21868_/B VGND VGND VPWR VPWR _22199_/X sky130_fd_sc_hd__or2_4
XFILLER_239_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16760_ _15061_/Y _16758_/X _16412_/X _16758_/X VGND VGND VPWR VPWR _24471_/D sky130_fd_sc_hd__a2bb2o_4
X_13972_ _14259_/A _13979_/D VGND VGND VPWR VPWR _15438_/C sky130_fd_sc_hd__or2_4
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20349__A3 _11851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15711_ _15710_/X VGND VGND VPWR VPWR _15854_/B sky130_fd_sc_hd__buf_2
X_12923_ _12787_/Y _12927_/B _12922_/Y VGND VGND VPWR VPWR _12923_/X sky130_fd_sc_hd__o21a_4
X_24909_ _24020_/CLK _24909_/D HRESETn VGND VGND VPWR VPWR _15618_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16691_ _24499_/Q VGND VGND VPWR VPWR _16691_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18430_ _18403_/X _18430_/B _18420_/X _18430_/D VGND VGND VPWR VPWR _18430_/X sky130_fd_sc_hd__or4_4
XANTENNA__25392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15642_ _21757_/A _15635_/X _15483_/X _15641_/X VGND VGND VPWR VPWR _15642_/X sky130_fd_sc_hd__a2bb2o_4
X_12854_ _12837_/Y _12796_/Y _12853_/Y VGND VGND VPWR VPWR _12854_/X sky130_fd_sc_hd__or3_4
XPHY_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14433__B1 _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15776__A3 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ HWDATA[16] VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__buf_2
X_18361_ _18361_/A _17491_/X VGND VGND VPWR VPWR _18361_/X sky130_fd_sc_hd__or2_4
XPHY_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15568_/Y _15572_/X _11755_/X _15572_/X VGND VGND VPWR VPWR _24928_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _25380_/Q _22428_/A _12783_/Y _12784_/Y VGND VGND VPWR VPWR _12785_/X sky130_fd_sc_hd__o22a_4
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19372__B1 _19305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17265_/X _17276_/X _17231_/Y VGND VGND VPWR VPWR _17313_/C sky130_fd_sc_hd__o21a_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14524_/A _14523_/X VGND VGND VPWR VPWR _25115_/D sky130_fd_sc_hd__or2_4
X_11736_ _11736_/A _11736_/B _11736_/C VGND VGND VPWR VPWR _11740_/C sky130_fd_sc_hd__or3_4
X_18292_ _18288_/X _17735_/X _18285_/D _17713_/X VGND VGND VPWR VPWR _24223_/D sky130_fd_sc_hd__o22a_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17227_/Y VGND VGND VPWR VPWR _17243_/X sky130_fd_sc_hd__buf_2
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _14455_/A VGND VGND VPWR VPWR _14455_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11667_ _13693_/A _24235_/Q _11666_/Y _24242_/Q VGND VGND VPWR VPWR _11675_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19124__B1 _19008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12747__B1 _12657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13332_/X _13402_/X _13406_/C VGND VGND VPWR VPWR _13406_/X sky130_fd_sc_hd__or3_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17173_/X VGND VGND VPWR VPWR _24378_/D sky130_fd_sc_hd__inv_2
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _14386_/A _21348_/A VGND VGND VPWR VPWR _14386_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_227_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _24337_/CLK sky130_fd_sc_hd__clkbuf_1
X_16125_ _24706_/Q VGND VGND VPWR VPWR _16125_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13337_ _13155_/X VGND VGND VPWR VPWR _13371_/A sky130_fd_sc_hd__buf_2
XFILLER_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12951__A _12828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16056_ _16044_/A VGND VGND VPWR VPWR _16056_/X sky130_fd_sc_hd__buf_2
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13207_/X _13266_/X _25337_/Q _13267_/X VGND VGND VPWR VPWR _13268_/X sky130_fd_sc_hd__o22a_4
X_15007_ _15256_/A _24451_/Q _15256_/A _24451_/Q VGND VGND VPWR VPWR _15011_/B sky130_fd_sc_hd__a2bb2o_4
X_12219_ _22418_/A VGND VGND VPWR VPWR _12219_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21234__B2 _15674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19734__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _13199_/A _23524_/Q VGND VGND VPWR VPWR _13199_/X sky130_fd_sc_hd__or2_4
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19815_ _19815_/A VGND VGND VPWR VPWR _19816_/A sky130_fd_sc_hd__inv_2
XFILLER_243_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13782__A _13782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17254__A _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16958_ _23237_/A _16957_/X _16166_/Y _24267_/Q VGND VGND VPWR VPWR _16958_/X sky130_fd_sc_hd__a2bb2o_4
X_19746_ _19745_/Y _19743_/X _19656_/X _19743_/X VGND VGND VPWR VPWR _23643_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15909_ _12778_/Y _15904_/X _15767_/X _15908_/X VGND VGND VPWR VPWR _24798_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19677_ _19032_/A VGND VGND VPWR VPWR _19677_/X sky130_fd_sc_hd__buf_2
X_16889_ _14791_/X VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__buf_2
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18628_ _24155_/Q VGND VGND VPWR VPWR _18682_/A sky130_fd_sc_hd__inv_2
XFILLER_80_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14424__B1 _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21504__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18559_ _18559_/A VGND VGND VPWR VPWR _18560_/B sky130_fd_sc_hd__inv_2
XANTENNA__19363__B1 _19341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21570_ _21570_/A VGND VGND VPWR VPWR _21570_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_37_0_HCLK clkbuf_6_36_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20521_ _24088_/Q _20520_/Y VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__and2_4
XFILLER_193_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17541__A1_N _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23240_ _23299_/A _23230_/X _23240_/C _23239_/X VGND VGND VPWR VPWR _23240_/X sky130_fd_sc_hd__or4_4
XFILLER_193_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20452_ _20444_/A _20451_/X VGND VGND VPWR VPWR _20455_/B sky130_fd_sc_hd__and2_4
XFILLER_119_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21877__C _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23171_ _22993_/X _23170_/X _23062_/X _11768_/A _23129_/X VGND VGND VPWR VPWR _23171_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_192_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20383_ _20383_/A VGND VGND VPWR VPWR _22364_/B sky130_fd_sc_hd__inv_2
XANTENNA__22670__B1 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22122_ _12952_/C _21027_/X _20855_/Y _22121_/X VGND VGND VPWR VPWR _22122_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22053_ _21526_/X _22053_/B VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__and2_4
XFILLER_88_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22422__B1 _22836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21004_ _21004_/A _14205_/X VGND VGND VPWR VPWR _23977_/D sky130_fd_sc_hd__and2_4
XFILLER_99_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16101__B1 _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22955_ _24540_/Q _22411_/X _15676_/X _22954_/X VGND VGND VPWR VPWR _22956_/C sky130_fd_sc_hd__a211o_4
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21906_ _22094_/A _21906_/B VGND VGND VPWR VPWR _21907_/C sky130_fd_sc_hd__or2_4
XFILLER_243_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22886_ _22436_/X _22874_/X _22886_/C _22885_/X VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__or4_4
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_238_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24625_ _24625_/CLK _16355_/X HRESETn VGND VGND VPWR VPWR _24625_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21837_ _13826_/X _21836_/X _24234_/Q _13824_/X VGND VGND VPWR VPWR _21838_/B sky130_fd_sc_hd__o22a_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19354__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12570_ _12583_/A _12568_/Y _12713_/A _12572_/A VGND VGND VPWR VPWR _12570_/X sky130_fd_sc_hd__a2bb2o_4
X_21768_ _21646_/A _21766_/X _21767_/X VGND VGND VPWR VPWR _21768_/X sky130_fd_sc_hd__and3_4
X_24556_ _24556_/CLK _24556_/D HRESETn VGND VGND VPWR VPWR _24556_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16168__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20719_ _15634_/Y _20716_/X _20704_/X _20718_/X VGND VGND VPWR VPWR _20720_/A sky130_fd_sc_hd__o22a_4
X_23507_ _24684_/CLK _20132_/X VGND VGND VPWR VPWR _20131_/A sky130_fd_sc_hd__dfxtp_4
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15915__B1 _21712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24785__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21699_ _22274_/A _21690_/X _21698_/X VGND VGND VPWR VPWR _21699_/X sky130_fd_sc_hd__or3_4
X_24487_ _24666_/CLK _24487_/D HRESETn VGND VGND VPWR VPWR _16720_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_211_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _25203_/Q VGND VGND VPWR VPWR _14240_/Y sky130_fd_sc_hd__inv_2
X_23438_ _23582_/CLK _23438_/D VGND VGND VPWR VPWR _20314_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24714__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14171_ _25219_/Q _14108_/B _25219_/Q _14108_/B VGND VGND VPWR VPWR _14171_/X sky130_fd_sc_hd__a2bb2o_4
X_23369_ VGND VGND VPWR VPWR _23369_/HI scl_o_S5 sky130_fd_sc_hd__conb_1
XFILLER_180_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_0_0_HCLK_A clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13122_ _13115_/B VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__inv_2
X_25108_ _23970_/CLK _14540_/X HRESETn VGND VGND VPWR VPWR _21352_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15143__B2 _16430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16340__B1 _16241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_57_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _24240_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_127_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13053_ _12998_/X _13061_/B VGND VGND VPWR VPWR _13053_/X sky130_fd_sc_hd__or2_4
X_17930_ _17930_/A _17929_/Y _17924_/B VGND VGND VPWR VPWR _17930_/X sky130_fd_sc_hd__or3_4
X_25039_ _25030_/CLK _25039_/D HRESETn VGND VGND VPWR VPWR _14910_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12004_ _12003_/X VGND VGND VPWR VPWR _12004_/Y sky130_fd_sc_hd__inv_2
X_17861_ _17861_/A _17861_/B _17861_/C _17861_/D VGND VGND VPWR VPWR _17864_/B sky130_fd_sc_hd__or4_4
XFILLER_239_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24957__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16812_ _14939_/Y _16806_/X HWDATA[29] _16811_/X VGND VGND VPWR VPWR _16812_/X sky130_fd_sc_hd__a2bb2o_4
X_19600_ _19599_/X VGND VGND VPWR VPWR _19615_/A sky130_fd_sc_hd__buf_2
XANTENNA__17074__A _17074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17792_ _17791_/X VGND VGND VPWR VPWR _17792_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19531_ _23715_/Q VGND VGND VPWR VPWR _22245_/B sky130_fd_sc_hd__inv_2
X_16743_ _16762_/A VGND VGND VPWR VPWR _16743_/X sky130_fd_sc_hd__buf_2
XFILLER_235_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13955_ _13955_/A _13955_/B _13954_/X _13962_/C VGND VGND VPWR VPWR _13955_/X sky130_fd_sc_hd__or4_4
XFILLER_207_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _12906_/A _12906_/B _12905_/X VGND VGND VPWR VPWR _25396_/D sky130_fd_sc_hd__and3_4
X_19462_ _19458_/Y _19461_/X _19439_/X _19461_/X VGND VGND VPWR VPWR _23740_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17802__A _16952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16674_ _16671_/Y _16667_/X _16315_/X _16673_/X VGND VGND VPWR VPWR _16674_/X sky130_fd_sc_hd__a2bb2o_4
X_13886_ _13880_/X _13885_/X _14277_/A _13876_/X VGND VGND VPWR VPWR _13886_/X sky130_fd_sc_hd__o22a_4
X_18413_ _16226_/A _24182_/Q _16226_/Y _18471_/A VGND VGND VPWR VPWR _18420_/A sky130_fd_sc_hd__o22a_4
X_15625_ _15625_/A VGND VGND VPWR VPWR _15625_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21324__A _21064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12837_ _25376_/Q VGND VGND VPWR VPWR _12837_/Y sky130_fd_sc_hd__inv_2
X_19393_ _19389_/Y _19392_/X _19326_/X _19392_/X VGND VGND VPWR VPWR _19393_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22139__B _21719_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11850__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18344_ _18333_/C _18333_/B _18959_/B VGND VGND VPWR VPWR _24212_/D sky130_fd_sc_hd__o21a_4
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15556_ _22891_/B VGND VGND VPWR VPWR _15758_/A sky130_fd_sc_hd__buf_2
X_12768_ _23199_/A VGND VGND VPWR VPWR _12768_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21152__B1 _25175_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14506_/X VGND VGND VPWR VPWR _14507_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11719_ _13607_/A VGND VGND VPWR VPWR _14199_/A sky130_fd_sc_hd__buf_2
X_18275_ _13804_/D _18262_/X _14248_/A _21514_/A _18269_/X VGND VGND VPWR VPWR _24227_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15906__B1 _15905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15487_ _14877_/Y _15485_/X _15486_/X _15485_/X VGND VGND VPWR VPWR _15487_/X sky130_fd_sc_hd__a2bb2o_4
X_12699_ _12618_/D _12674_/X _12657_/A _12697_/B VGND VGND VPWR VPWR _12700_/A sky130_fd_sc_hd__a211o_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17226_ _16317_/Y _17231_/A _16348_/A _17359_/C VGND VGND VPWR VPWR _17226_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14438_ _14437_/Y _14435_/X _14248_/X _14435_/X VGND VGND VPWR VPWR _25144_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22155__A _24622_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17157_ _17157_/A _17155_/Y _17160_/C VGND VGND VPWR VPWR _24384_/D sky130_fd_sc_hd__and3_4
X_14369_ _14369_/A VGND VGND VPWR VPWR _14369_/X sky130_fd_sc_hd__buf_2
XFILLER_155_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16153__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16108_ _23205_/A VGND VGND VPWR VPWR _16108_/Y sky130_fd_sc_hd__inv_2
X_17088_ _17088_/A _17088_/B VGND VGND VPWR VPWR _17088_/X sky130_fd_sc_hd__or2_4
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15685__A2 _15678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16039_ _16038_/Y _16036_/X _15970_/X _16036_/X VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16882__B2 _16877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22955__A1 _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19729_ _19727_/Y _19725_/X _19728_/X _19725_/X VGND VGND VPWR VPWR _19729_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17712__A _17712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22740_ _24600_/Q _22827_/B VGND VGND VPWR VPWR _22743_/B sky130_fd_sc_hd__or2_4
XFILLER_92_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22671_ _22671_/A VGND VGND VPWR VPWR _22671_/Y sky130_fd_sc_hd__inv_2
XFILLER_240_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18854__A1_N _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19336__B1 _19246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21622_ _21648_/A _21622_/B VGND VGND VPWR VPWR _21622_/X sky130_fd_sc_hd__or2_4
X_24410_ _24642_/CLK _24410_/D HRESETn VGND VGND VPWR VPWR _21022_/B sky130_fd_sc_hd__dfrtp_4
X_25390_ _25392_/CLK _25390_/D HRESETn VGND VGND VPWR VPWR _12819_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21553_ _21542_/X _21546_/Y _22723_/A _21552_/X VGND VGND VPWR VPWR _21553_/X sky130_fd_sc_hd__a2bb2o_4
X_24341_ _24343_/CLK _17418_/X HRESETn VGND VGND VPWR VPWR _24341_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__19639__A _19639_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20504_ _20504_/A _20494_/Y _24088_/Q VGND VGND VPWR VPWR _20505_/B sky130_fd_sc_hd__and3_4
X_24272_ _24272_/CLK _24272_/D HRESETn VGND VGND VPWR VPWR _17871_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21484_ _21676_/A _19960_/Y VGND VGND VPWR VPWR _21484_/X sky130_fd_sc_hd__or2_4
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16570__B1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23223_ _24478_/Q _23016_/X _23190_/X VGND VGND VPWR VPWR _23223_/X sky130_fd_sc_hd__o21a_4
X_20435_ _20434_/Y _20430_/X _20249_/X _20430_/A VGND VGND VPWR VPWR _20435_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_210_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24566_/CLK sky130_fd_sc_hd__clkbuf_1
X_23154_ _24444_/Q _22947_/X _23015_/X _23153_/X VGND VGND VPWR VPWR _23154_/X sky130_fd_sc_hd__a211o_4
X_20366_ _20362_/Y _20365_/X _19626_/A _20365_/X VGND VGND VPWR VPWR _20366_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22105_ _21879_/A _22102_/X _22105_/C VGND VGND VPWR VPWR _22105_/X sky130_fd_sc_hd__and3_4
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23085_ _23065_/X _23068_/X _23072_/Y _23084_/X VGND VGND VPWR VPWR HRDATA[23] sky130_fd_sc_hd__a211o_4
X_20297_ _14804_/Y _23985_/Q VGND VGND VPWR VPWR _20297_/X sky130_fd_sc_hd__or2_4
X_22036_ _22036_/A _22036_/B _22036_/C VGND VGND VPWR VPWR _22036_/X sky130_fd_sc_hd__and3_4
XFILLER_102_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19811__B2 _19806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11935__A _11934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15979__A3 _16241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23987_ _23991_/CLK _20626_/Y HRESETn VGND VGND VPWR VPWR _20624_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22174__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ _11691_/A _13740_/B VGND VGND VPWR VPWR _13740_/X sky130_fd_sc_hd__or2_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15143__A2_N _16430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22938_ _23008_/A _22938_/B VGND VGND VPWR VPWR _22938_/Y sky130_fd_sc_hd__nor2_4
XFILLER_216_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20185__B2 _20184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13671_ _13671_/A _13671_/B VGND VGND VPWR VPWR _13671_/X sky130_fd_sc_hd__or2_4
XFILLER_204_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22869_ _22860_/Y _22867_/Y _22868_/X VGND VGND VPWR VPWR _22869_/X sky130_fd_sc_hd__o21a_4
XFILLER_232_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16238__A _16238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19327__B1 _19326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15410_ _15393_/A _15407_/B _15409_/Y VGND VGND VPWR VPWR _24990_/D sky130_fd_sc_hd__and3_4
X_12622_ _12622_/A VGND VGND VPWR VPWR _12623_/D sky130_fd_sc_hd__inv_2
X_24608_ _24602_/CLK _24608_/D HRESETn VGND VGND VPWR VPWR _24608_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16390_ _16390_/A VGND VGND VPWR VPWR _16415_/A sky130_fd_sc_hd__buf_2
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15341_ _15355_/A _15341_/B _15340_/X VGND VGND VPWR VPWR _15341_/X sky130_fd_sc_hd__and3_4
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17889__B1 _16964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12553_ _12543_/X _12553_/B _12549_/X _12553_/D VGND VGND VPWR VPWR _12553_/X sky130_fd_sc_hd__or4_4
X_24539_ _24537_/CLK _16585_/X HRESETn VGND VGND VPWR VPWR _24539_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18060_ _18060_/A _19150_/A VGND VGND VPWR VPWR _18060_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_20_0_HCLK clkbuf_5_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _15255_/X _15270_/X _15271_/X VGND VGND VPWR VPWR _25022_/D sky130_fd_sc_hd__and3_4
XFILLER_8_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12287_/A _12481_/X VGND VGND VPWR VPWR _12485_/C sky130_fd_sc_hd__or2_4
XANTENNA__16561__B1 _16389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__A1 _12132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15903__A3 _16252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17011_ _16046_/Y _24393_/Q _16046_/Y _24393_/Q VGND VGND VPWR VPWR _17011_/X sky130_fd_sc_hd__a2bb2o_4
X_14223_ _14223_/A VGND VGND VPWR VPWR _21004_/A sky130_fd_sc_hd__inv_2
XFILLER_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14154_ _14134_/X _14152_/Y _14111_/A _14153_/X VGND VGND VPWR VPWR _14154_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16313__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13105_ _12332_/Y _13092_/X VGND VGND VPWR VPWR _13105_/Y sky130_fd_sc_hd__nand2_4
X_14085_ _14069_/B VGND VGND VPWR VPWR _14085_/X sky130_fd_sc_hd__buf_2
X_18962_ _18958_/Y _18961_/X _17427_/X _18961_/X VGND VGND VPWR VPWR _18962_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_152_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22937__B2 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13036_ _13036_/A VGND VGND VPWR VPWR _25366_/D sky130_fd_sc_hd__inv_2
X_17913_ _17910_/B _17913_/B VGND VGND VPWR VPWR _17915_/A sky130_fd_sc_hd__or2_4
X_18893_ _18893_/A VGND VGND VPWR VPWR _18893_/X sky130_fd_sc_hd__buf_2
X_17844_ _17852_/A _17844_/B _17844_/C VGND VGND VPWR VPWR _24278_/D sky130_fd_sc_hd__and3_4
XFILLER_227_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16092__A2 _21596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17775_ _16925_/Y _16957_/X _17775_/C _17774_/X VGND VGND VPWR VPWR _17776_/A sky130_fd_sc_hd__or4_4
X_14987_ _14986_/Y _24449_/Q _14986_/Y _24449_/Q VGND VGND VPWR VPWR _14987_/X sky130_fd_sc_hd__a2bb2o_4
X_16726_ _14479_/A VGND VGND VPWR VPWR _16726_/X sky130_fd_sc_hd__buf_2
X_19514_ _22022_/B _19508_/X _11948_/X _19513_/X VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13938_ _13967_/C VGND VGND VPWR VPWR _13948_/C sky130_fd_sc_hd__buf_2
XFILLER_241_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19445_ _19443_/Y _19438_/X _19421_/X _19444_/X VGND VGND VPWR VPWR _19445_/X sky130_fd_sc_hd__a2bb2o_4
X_16657_ _24513_/Q VGND VGND VPWR VPWR _16657_/Y sky130_fd_sc_hd__inv_2
X_13869_ _24008_/Q VGND VGND VPWR VPWR _13869_/X sky130_fd_sc_hd__buf_2
XFILLER_234_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_205_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15608_ _15608_/A VGND VGND VPWR VPWR _15608_/Y sky130_fd_sc_hd__inv_2
X_19376_ _19376_/A VGND VGND VPWR VPWR _19376_/Y sky130_fd_sc_hd__inv_2
X_16588_ _24537_/Q VGND VGND VPWR VPWR _16588_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24636__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18327_ _18326_/X VGND VGND VPWR VPWR _18327_/Y sky130_fd_sc_hd__inv_2
X_15539_ _15537_/Y _15533_/X HADDR[7] _15538_/X VGND VGND VPWR VPWR _15539_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20182__A2_N _20177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22873__B1 _24843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _18241_/Y VGND VGND VPWR VPWR _18258_/X sky130_fd_sc_hd__buf_2
XFILLER_175_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17209_ _24619_/Q _24348_/Q _16370_/Y _17389_/A VGND VGND VPWR VPWR _17210_/D sky130_fd_sc_hd__o22a_4
X_18189_ _18189_/A _18189_/B VGND VGND VPWR VPWR _18191_/B sky130_fd_sc_hd__or2_4
X_20220_ _20218_/Y _20214_/X _16874_/X _20219_/X VGND VGND VPWR VPWR _23474_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20151_ _20150_/Y VGND VGND VPWR VPWR _20151_/X sky130_fd_sc_hd__buf_2
XANTENNA__25495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22410__A1_N _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_40_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23475_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20082_ _20078_/Y _20081_/X _19817_/X _20081_/X VGND VGND VPWR VPWR _23524_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20120__A2_N _20118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23050__B1 _24848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23910_ _24111_/CLK _18978_/X VGND VGND VPWR VPWR _23910_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11755__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24890_ _24872_/CLK _15724_/X HRESETn VGND VGND VPWR VPWR _24890_/Q sky130_fd_sc_hd__dfrtp_4
X_23841_ _24100_/CLK _19177_/X VGND VGND VPWR VPWR _18100_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20984_ _12164_/X _20982_/B VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__and2_4
X_23772_ _25077_/CLK _19370_/X VGND VGND VPWR VPWR _17955_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21364__B1 _12175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25511_ _23408_/CLK _25511_/D HRESETn VGND VGND VPWR VPWR _20003_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22723_ _22723_/A _22723_/B _22722_/X VGND VGND VPWR VPWR _22723_/X sky130_fd_sc_hd__and3_4
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11852__B1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16058__A _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25442_ _25444_/CLK _12506_/Y HRESETn VGND VGND VPWR VPWR _25442_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21899__A _22093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22654_ _22768_/A _22654_/B VGND VGND VPWR VPWR _22654_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21605_ _21605_/A VGND VGND VPWR VPWR _21605_/X sky130_fd_sc_hd__buf_2
XFILLER_185_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22585_ _12855_/C _22678_/B _22584_/X VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__o21a_4
X_25373_ _24799_/CLK _25373_/D HRESETn VGND VGND VPWR VPWR _21035_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24324_ _23534_/CLK _17613_/Y HRESETn VGND VGND VPWR VPWR _24324_/Q sky130_fd_sc_hd__dfrtp_4
X_21536_ _21543_/A VGND VGND VPWR VPWR _21536_/X sky130_fd_sc_hd__buf_2
XANTENNA__16543__B1 _16368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21467_ _21466_/X _21467_/B VGND VGND VPWR VPWR _21467_/X sky130_fd_sc_hd__or2_4
X_24255_ _24258_/CLK _17937_/X HRESETn VGND VGND VPWR VPWR _17929_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_181_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20418_ _20408_/X _21382_/B _13481_/A _21218_/A _20406_/A VGND VGND VPWR VPWR _20418_/X
+ sky130_fd_sc_hd__a32o_4
X_23206_ _22993_/X _23205_/X _23062_/X _25552_/Q _23129_/X VGND VGND VPWR VPWR _23206_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21398_ _21240_/A VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__buf_2
X_24186_ _23973_/CLK _18524_/X HRESETn VGND VGND VPWR VPWR _24186_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12580__B2 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20349_ _20342_/X _19599_/D _11851_/A _21996_/C _20346_/X VGND VGND VPWR VPWR _23425_/D
+ sky130_fd_sc_hd__a32o_4
X_23137_ _22476_/A VGND VGND VPWR VPWR _23137_/X sky130_fd_sc_hd__buf_2
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23068_ _23066_/X _23068_/B _22929_/X VGND VGND VPWR VPWR _23068_/X sky130_fd_sc_hd__or3_4
XANTENNA__23041__B1 _12377_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14910_ _14910_/A VGND VGND VPWR VPWR _14910_/Y sky130_fd_sc_hd__inv_2
X_22019_ _21212_/A VGND VGND VPWR VPWR _22265_/A sky130_fd_sc_hd__buf_2
XFILLER_248_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19832__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15890_ _15880_/A VGND VGND VPWR VPWR _15890_/X sky130_fd_sc_hd__buf_2
X_14841_ _14812_/C _14826_/X _14828_/A _14827_/Y VGND VGND VPWR VPWR _14841_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13880__A _24007_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17560_ _17560_/A _17560_/B _17558_/X _17560_/D VGND VGND VPWR VPWR _17561_/D sky130_fd_sc_hd__or4_4
XFILLER_17_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12096__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14772_ _14772_/A _14781_/A _14772_/C VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__or3_4
X_11984_ _11970_/C _11979_/C _11984_/C VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__or3_4
XFILLER_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16511_ _16510_/Y _16508_/X _16238_/X _16508_/X VGND VGND VPWR VPWR _24567_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ _13722_/X VGND VGND VPWR VPWR _13723_/X sky130_fd_sc_hd__buf_2
X_17491_ _17485_/Y _17459_/A _11658_/A VGND VGND VPWR VPWR _17491_/X sky130_fd_sc_hd__and3_4
XANTENNA__11843__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19230_ _19230_/A VGND VGND VPWR VPWR _19230_/Y sky130_fd_sc_hd__inv_2
X_16442_ _16442_/A VGND VGND VPWR VPWR _16442_/X sky130_fd_sc_hd__buf_2
X_13654_ _25303_/Q _13533_/X _13649_/X VGND VGND VPWR VPWR _13654_/X sky130_fd_sc_hd__a21o_4
XFILLER_177_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12605_ _12599_/Y VGND VGND VPWR VPWR _12740_/A sky130_fd_sc_hd__buf_2
X_19161_ _19161_/A VGND VGND VPWR VPWR _19161_/Y sky130_fd_sc_hd__inv_2
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _16372_/Y _16291_/A _16276_/X _16291_/A VGND VGND VPWR VPWR _24618_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22855__B1 _22852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13585_ _25096_/Q VGND VGND VPWR VPWR _14603_/A sky130_fd_sc_hd__inv_2
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18183__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18112_ _18037_/A _18112_/B _18112_/C VGND VGND VPWR VPWR _18112_/X sky130_fd_sc_hd__and3_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15324_ _15357_/A VGND VGND VPWR VPWR _15324_/X sky130_fd_sc_hd__buf_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12536_ _12536_/A VGND VGND VPWR VPWR _12536_/Y sky130_fd_sc_hd__inv_2
X_19092_ _19089_/Y _19090_/X _19091_/X _19090_/X VGND VGND VPWR VPWR _19092_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18043_ _18209_/A _23754_/Q VGND VGND VPWR VPWR _18043_/X sky130_fd_sc_hd__or2_4
X_15255_ _15293_/A VGND VGND VPWR VPWR _15255_/X sky130_fd_sc_hd__buf_2
X_12467_ _12467_/A VGND VGND VPWR VPWR _12467_/Y sky130_fd_sc_hd__inv_2
X_14206_ _20675_/A VGND VGND VPWR VPWR _14816_/A sky130_fd_sc_hd__inv_2
X_15186_ _15182_/B _15174_/X VGND VGND VPWR VPWR _15186_/X sky130_fd_sc_hd__or2_4
XFILLER_153_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12398_ _12398_/A _12398_/B _12398_/C VGND VGND VPWR VPWR _25469_/D sky130_fd_sc_hd__and3_4
XFILLER_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20094__B1 _19734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14137_ _25149_/Q VGND VGND VPWR VPWR _14137_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19994_ _22256_/B _19989_/X _19993_/X _19989_/X VGND VGND VPWR VPWR _23555_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_27_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14068_ _14068_/A VGND VGND VPWR VPWR _14069_/B sky130_fd_sc_hd__buf_2
X_18945_ _18952_/A VGND VGND VPWR VPWR _18945_/X sky130_fd_sc_hd__buf_2
X_13019_ _13019_/A _13013_/B _13019_/C VGND VGND VPWR VPWR _13020_/A sky130_fd_sc_hd__or3_4
XFILLER_228_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21991__B _21991_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18876_ _18876_/A VGND VGND VPWR VPWR _18876_/X sky130_fd_sc_hd__buf_2
XFILLER_95_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21594__B1 _21591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17827_ _17827_/A VGND VGND VPWR VPWR _17827_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24888__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15273__B1 _14996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17758_ _24266_/Q VGND VGND VPWR VPWR _17758_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21346__B1 _15676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24817__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16709_ _16709_/A VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__buf_2
X_17689_ _17687_/A _17676_/X _17689_/C VGND VGND VPWR VPWR _17689_/X sky130_fd_sc_hd__and3_4
XFILLER_23_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15025__B1 _15292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19428_ _18149_/B VGND VGND VPWR VPWR _19428_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19359_ _23775_/Q VGND VGND VPWR VPWR _19359_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22310__A2 _22301_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16606__A _16606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22370_ _17738_/A _22349_/Y _22356_/Y _22363_/Y _22369_/Y VGND VGND VPWR VPWR _22370_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21321_ _21321_/A VGND VGND VPWR VPWR _21321_/X sky130_fd_sc_hd__buf_2
XFILLER_163_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21252_ _21244_/X _21250_/X _21251_/X VGND VGND VPWR VPWR _21252_/X sky130_fd_sc_hd__o21a_4
X_24040_ _24042_/CLK _20807_/X HRESETn VGND VGND VPWR VPWR _13145_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20203_ _21783_/B _20198_/X _20115_/X _20198_/X VGND VGND VPWR VPWR _23480_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12248__A1_N _12247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21183_ _17714_/A _21181_/X _21183_/C VGND VGND VPWR VPWR _21183_/X sky130_fd_sc_hd__and3_4
XANTENNA__16341__A _24630_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22062__B _23354_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20134_ _20129_/A VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__buf_2
XANTENNA__19778__B1 _19753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13511__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20065_ _20059_/Y VGND VGND VPWR VPWR _20065_/X sky130_fd_sc_hd__buf_2
X_24942_ _23408_/CLK _15527_/X HRESETn VGND VGND VPWR VPWR _15524_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_219_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24873_ _24872_/CLK _15757_/X HRESETn VGND VGND VPWR VPWR _24873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14796__A _18059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15803__A2 _15797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23824_ _23830_/CLK _23824_/D VGND VGND VPWR VPWR _18136_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24558__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21337__B1 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23669_/CLK _23755_/D VGND VGND VPWR VPWR _23755_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20836_/X _20966_/X _16651_/A _20883_/A VGND VGND VPWR VPWR _24077_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12816__A1_N _22678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22706_ _13571_/Y _22706_/B VGND VGND VPWR VPWR _22706_/X sky130_fd_sc_hd__and2_4
XANTENNA__15567__A1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ _23703_/CLK _23686_/D VGND VGND VPWR VPWR _19617_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_202_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20895_/Y _20896_/Y _20897_/X VGND VGND VPWR VPWR _20898_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22518__A _16284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25425_ _25425_/CLK _12687_/X HRESETn VGND VGND VPWR VPWR _12541_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21422__A _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22637_ _24664_/Q _22589_/B VGND VGND VPWR VPWR _22640_/B sky130_fd_sc_hd__or2_4
XFILLER_213_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13370_ _13254_/X _13368_/X _13370_/C VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__and3_4
X_25356_ _25358_/CLK _13073_/X HRESETn VGND VGND VPWR VPWR _25356_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16516__B1 _16245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22568_ _22568_/A _21450_/X VGND VGND VPWR VPWR _22568_/X sky130_fd_sc_hd__or2_4
XFILLER_210_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12321_ _13088_/A _24825_/Q _13088_/A _24825_/Q VGND VGND VPWR VPWR _12321_/X sky130_fd_sc_hd__a2bb2o_4
X_24307_ _24302_/CLK _17681_/X HRESETn VGND VGND VPWR VPWR _24307_/Q sky130_fd_sc_hd__dfrtp_4
X_21519_ _21180_/X VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__buf_2
X_25287_ _24233_/CLK _25287_/D HRESETn VGND VGND VPWR VPWR _11691_/A sky130_fd_sc_hd__dfrtp_4
X_22499_ _22494_/X _22496_/X _22497_/X _24730_/Q _22498_/X VGND VGND VPWR VPWR _22500_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_6_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20980__B _12168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15040_ _25023_/Q VGND VGND VPWR VPWR _15260_/C sky130_fd_sc_hd__inv_2
XFILLER_108_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12252_ _12439_/A _22665_/A _12439_/A _22665_/A VGND VGND VPWR VPWR _12260_/A sky130_fd_sc_hd__a2bb2o_4
X_24238_ _24238_/CLK _24238_/D HRESETn VGND VGND VPWR VPWR _24238_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12183_ SSn_S3 _12182_/Y _11871_/X _12182_/Y VGND VGND VPWR VPWR _12183_/X sky130_fd_sc_hd__a2bb2o_4
X_24169_ _24169_/CLK _18586_/X HRESETn VGND VGND VPWR VPWR _24169_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16991_ _16010_/A _16990_/A _16010_/Y _17072_/A VGND VGND VPWR VPWR _16998_/A sky130_fd_sc_hd__o22a_4
X_15942_ _15938_/X _15902_/X _15562_/X _24784_/Q _15941_/X VGND VGND VPWR VPWR _24784_/D
+ sky130_fd_sc_hd__a32o_4
X_18730_ _18701_/X _18710_/X _18702_/A VGND VGND VPWR VPWR _18731_/C sky130_fd_sc_hd__o21a_4
XFILLER_89_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18661_ _24159_/Q VGND VGND VPWR VPWR _18670_/A sky130_fd_sc_hd__inv_2
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18441__B1 _24673_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15873_ _15858_/X _15865_/X _15562_/X _24821_/Q _15872_/X VGND VGND VPWR VPWR _24821_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14824_ _14824_/A _14824_/B _25054_/Q VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__or3_4
X_17612_ _17569_/A _17610_/X _17611_/X _17606_/B VGND VGND VPWR VPWR _17613_/A sky130_fd_sc_hd__a211o_4
X_18592_ _18433_/Y _18565_/X VGND VGND VPWR VPWR _18597_/B sky130_fd_sc_hd__or2_4
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24910__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17543_ _11816_/Y _17666_/A _11816_/Y _17666_/A VGND VGND VPWR VPWR _17547_/A sky130_fd_sc_hd__a2bb2o_4
X_14755_ _14693_/Y _14755_/B VGND VGND VPWR VPWR _14755_/X sky130_fd_sc_hd__or2_4
XFILLER_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11967_ _11967_/A VGND VGND VPWR VPWR _11979_/A sky130_fd_sc_hd__buf_2
XFILLER_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13706_ _13685_/Y _13689_/X _13703_/A _25301_/Q _13705_/Y VGND VGND VPWR VPWR _13706_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_232_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17474_ _13183_/X _17461_/X _18347_/A VGND VGND VPWR VPWR _17474_/X sky130_fd_sc_hd__o21a_4
XFILLER_205_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14686_ _14692_/A VGND VGND VPWR VPWR _14686_/X sky130_fd_sc_hd__buf_2
XANTENNA__16755__B1 _15738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11898_ _11898_/A _11898_/B VGND VGND VPWR VPWR _11898_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22428__A _22428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ _24600_/Q VGND VGND VPWR VPWR _16425_/Y sky130_fd_sc_hd__inv_2
X_19213_ _19209_/Y _19212_/X _19169_/X _19212_/X VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21332__A _21332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13637_ _25079_/Q VGND VGND VPWR VPWR _19143_/A sky130_fd_sc_hd__buf_2
X_19144_ _19143_/X VGND VGND VPWR VPWR _19159_/A sky130_fd_sc_hd__inv_2
X_16356_ _24624_/Q VGND VGND VPWR VPWR _16356_/Y sky130_fd_sc_hd__inv_2
X_13568_ _25093_/Q VGND VGND VPWR VPWR _14610_/A sky130_fd_sc_hd__inv_2
XFILLER_146_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15307_ _15365_/A _15362_/A _15306_/X VGND VGND VPWR VPWR _15307_/X sky130_fd_sc_hd__or3_4
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12519_ _12519_/A VGND VGND VPWR VPWR _12623_/C sky130_fd_sc_hd__inv_2
X_19075_ _18938_/A _19075_/B _18938_/C VGND VGND VPWR VPWR _19075_/X sky130_fd_sc_hd__or3_4
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16287_ _24648_/Q VGND VGND VPWR VPWR _16287_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13499_ _13497_/Y _13498_/X _11867_/X _13498_/X VGND VGND VPWR VPWR _25324_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18026_ _13625_/X _18023_/X _18026_/C VGND VGND VPWR VPWR _18026_/X sky130_fd_sc_hd__and3_4
X_15238_ _15231_/A _15219_/X _15208_/X _15235_/Y VGND VGND VPWR VPWR _15238_/X sky130_fd_sc_hd__a211o_4
XANTENNA__25087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13785__A _19550_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ _15415_/A _24591_/Q _15310_/A _24588_/Q VGND VGND VPWR VPWR _15169_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18275__A3 _14248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16161__A _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12600__A2_N _24863_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19977_ _19976_/Y _19972_/X _19639_/X _19972_/X VGND VGND VPWR VPWR _19977_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18928_ _23927_/Q VGND VGND VPWR VPWR _18928_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22610__B _22610_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21507__A _21815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18859_ _16529_/Y _24138_/Q _16529_/Y _24138_/Q VGND VGND VPWR VPWR _18861_/C sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_114_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24923_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_216_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_177_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _25181_/CLK sky130_fd_sc_hd__clkbuf_1
X_21870_ _21870_/A _21855_/B _21752_/B VGND VGND VPWR VPWR _21870_/X sky130_fd_sc_hd__and3_4
XFILLER_227_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24651__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20821_ _20822_/A VGND VGND VPWR VPWR _20821_/Y sky130_fd_sc_hd__inv_2
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23540_ _23563_/CLK _23540_/D VGND VGND VPWR VPWR _23540_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ _20752_/A VGND VGND VPWR VPWR _20752_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16746__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ _20683_/A _20683_/B _20682_/X VGND VGND VPWR VPWR _20683_/X sky130_fd_sc_hd__and3_4
X_23471_ _23799_/CLK _23471_/D VGND VGND VPWR VPWR _20225_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25210_ _25200_/CLK _14220_/X HRESETn VGND VGND VPWR VPWR _14218_/A sky130_fd_sc_hd__dfrtp_4
X_22422_ _21082_/X _22419_/X _22836_/A _22421_/X VGND VGND VPWR VPWR _22422_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25141_ _25148_/CLK _25141_/D HRESETn VGND VGND VPWR VPWR _25141_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_164_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22353_ _21947_/A _22353_/B VGND VGND VPWR VPWR _22353_/X sky130_fd_sc_hd__or2_4
XFILLER_109_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21304_ _21296_/X _21304_/B _21308_/C VGND VGND VPWR VPWR _21304_/X sky130_fd_sc_hd__and3_4
XFILLER_164_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22284_ _21450_/X VGND VGND VPWR VPWR _22284_/X sky130_fd_sc_hd__buf_2
X_25072_ _23703_/CLK _14748_/X HRESETn VGND VGND VPWR VPWR _14734_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15721__A1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23169__A _22155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22598__A2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21235_ _11744_/X VGND VGND VPWR VPWR _21235_/X sky130_fd_sc_hd__buf_2
X_24023_ _24493_/CLK _20734_/Y HRESETn VGND VGND VPWR VPWR _20730_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18266__A3 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21166_ _17447_/Y _21134_/Y _14199_/B _21165_/X VGND VGND VPWR VPWR _21177_/A sky130_fd_sc_hd__a211o_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22801__A _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20117_ _23511_/Q VGND VGND VPWR VPWR _20117_/Y sky130_fd_sc_hd__inv_2
XFILLER_219_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21097_ _21023_/A _21109_/B VGND VGND VPWR VPWR _21097_/X sky130_fd_sc_hd__and2_4
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24739__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_73_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20048_ _23536_/Q VGND VGND VPWR VPWR _21807_/B sky130_fd_sc_hd__inv_2
X_24925_ _24825_/CLK _24925_/D HRESETn VGND VGND VPWR VPWR _24925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_219_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17226__B2 _17359_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12870_ _12906_/A _12868_/X _12869_/X VGND VGND VPWR VPWR _12870_/X sky130_fd_sc_hd__and3_4
X_24856_ _24856_/CLK _24856_/D HRESETn VGND VGND VPWR VPWR _24856_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ HWDATA[12] VGND VGND VPWR VPWR _16248_/A sky130_fd_sc_hd__buf_2
X_23807_ _23799_/CLK _23807_/D VGND VGND VPWR VPWR _19270_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24787_/CLK _15932_/X HRESETn VGND VGND VPWR VPWR _21023_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _21526_/X _21998_/X _21520_/X VGND VGND VPWR VPWR _21999_/Y sky130_fd_sc_hd__a21oi_4
XPHY_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14530_/X _14539_/X _14499_/A _14515_/Y VGND VGND VPWR VPWR _14540_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ HWDATA[31] VGND VGND VPWR VPWR _11752_/X sky130_fd_sc_hd__buf_2
X_23738_ _23794_/CLK _23738_/D VGND VGND VPWR VPWR _18046_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14470_/Y _14468_/X _14400_/X _14468_/X VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11682_/Y _22707_/A _11682_/Y _22707_/A VGND VGND VPWR VPWR _11684_/D sky130_fd_sc_hd__a2bb2o_4
X_23669_ _23669_/CLK _23669_/D VGND VGND VPWR VPWR _13461_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16227_/A VGND VGND VPWR VPWR _16210_/X sky130_fd_sc_hd__buf_2
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13454_/A _13422_/B _13422_/C VGND VGND VPWR VPWR _13423_/C sky130_fd_sc_hd__and3_4
X_25408_ _25410_/CLK _12743_/X HRESETn VGND VGND VPWR VPWR _25408_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17190_ _17190_/A _17185_/X _17188_/X _17190_/D VGND VGND VPWR VPWR _17211_/B sky130_fd_sc_hd__or4_4
XANTENNA__25527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16141_ _16162_/A VGND VGND VPWR VPWR _16141_/X sky130_fd_sc_hd__buf_2
XFILLER_210_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13353_ _13385_/A _13353_/B VGND VGND VPWR VPWR _13353_/X sky130_fd_sc_hd__or2_4
X_25339_ _24029_/CLK _13151_/X HRESETn VGND VGND VPWR VPWR _21130_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _13014_/A _24856_/Q _13014_/A _24856_/Q VGND VGND VPWR VPWR _12310_/B sky130_fd_sc_hd__a2bb2o_4
X_16072_ _24726_/Q VGND VGND VPWR VPWR _16072_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13284_ _13391_/A _13284_/B _13283_/X VGND VGND VPWR VPWR _13285_/C sky130_fd_sc_hd__or3_4
X_15023_ _15270_/A _15022_/A _15271_/A _15022_/Y VGND VGND VPWR VPWR _15030_/A sky130_fd_sc_hd__o22a_4
X_19900_ _19900_/A VGND VGND VPWR VPWR _19900_/X sky130_fd_sc_hd__buf_2
X_12235_ _12224_/X _12235_/B _12231_/X _12235_/D VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__or4_4
XANTENNA__22414__C _22303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19831_ _23614_/Q VGND VGND VPWR VPWR _19831_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12166_ _12166_/A _12166_/B _24120_/D _12166_/D VGND VGND VPWR VPWR _14342_/B sky130_fd_sc_hd__or4_4
XANTENNA__17465__B2 _13186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19762_ _19760_/Y _19756_/X _19761_/X _19742_/Y VGND VGND VPWR VPWR _23637_/D sky130_fd_sc_hd__a2bb2o_4
X_12097_ _12097_/A VGND VGND VPWR VPWR _12097_/Y sky130_fd_sc_hd__inv_2
X_16974_ _16974_/A VGND VGND VPWR VPWR _17050_/D sky130_fd_sc_hd__inv_2
XFILLER_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25139__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18713_ _18713_/A VGND VGND VPWR VPWR _18714_/A sky130_fd_sc_hd__inv_2
XFILLER_237_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21327__A _16731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15925_ _15924_/X VGND VGND VPWR VPWR _15925_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19693_ _19691_/Y _19689_/X _19692_/X _19689_/X VGND VGND VPWR VPWR _23662_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22761__A2 _22760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _15683_/X _15854_/B VGND VGND VPWR VPWR _15856_/X sky130_fd_sc_hd__or2_4
X_18644_ _18768_/A VGND VGND VPWR VPWR _18764_/A sky130_fd_sc_hd__inv_2
XFILLER_76_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14807_ _14873_/A _14873_/B _14889_/A _25049_/Q VGND VGND VPWR VPWR _14822_/B sky130_fd_sc_hd__or4_4
XANTENNA__24062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _15561_/Y _15664_/X _15782_/X _23386_/D _15786_/X VGND VGND VPWR VPWR _24858_/D
+ sky130_fd_sc_hd__a32o_4
X_18575_ _18479_/C _18573_/X _18574_/Y VGND VGND VPWR VPWR _18575_/X sky130_fd_sc_hd__o21a_4
X_12999_ _12996_/Y _13054_/A _12998_/X VGND VGND VPWR VPWR _12999_/X sky130_fd_sc_hd__or3_4
X_14738_ _22056_/A _14749_/B VGND VGND VPWR VPWR _14738_/Y sky130_fd_sc_hd__nand2_4
X_17526_ _25554_/Q _17525_/A _11757_/Y _17525_/Y VGND VGND VPWR VPWR _17526_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23261__B _23087_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17457_ _13607_/A _21178_/A VGND VGND VPWR VPWR _17458_/C sky130_fd_sc_hd__or2_4
X_14669_ _13611_/A VGND VGND VPWR VPWR _19028_/B sky130_fd_sc_hd__buf_2
XFILLER_177_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16408_ _15158_/Y _16403_/X _16407_/X _16403_/X VGND VGND VPWR VPWR _24607_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17388_ _17253_/Y _17390_/B _17387_/Y VGND VGND VPWR VPWR _24349_/D sky130_fd_sc_hd__o21a_4
X_16339_ _16352_/A VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__buf_2
X_19127_ _19125_/Y _19121_/X _19012_/X _19126_/X VGND VGND VPWR VPWR _19127_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22605__B _21104_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19058_ _23883_/Q VGND VGND VPWR VPWR _19058_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ _18126_/A _23883_/Q VGND VGND VPWR VPWR _18010_/C sky130_fd_sc_hd__or2_4
XFILLER_160_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21020_ _21020_/A _21020_/B VGND VGND VPWR VPWR _21020_/X sky130_fd_sc_hd__and2_4
XANTENNA__18653__B1 _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17715__A _21212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24832__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22971_ _22837_/X _22962_/Y _22966_/Y _22970_/X VGND VGND VPWR VPWR _22979_/C sky130_fd_sc_hd__a211o_4
XFILLER_95_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24710_ _25444_/CLK _24710_/D HRESETn VGND VGND VPWR VPWR _24710_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11763__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21922_ _21895_/X _21922_/B VGND VGND VPWR VPWR _21922_/X sky130_fd_sc_hd__or2_4
XFILLER_83_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24641_ _24641_/CLK _24641_/D HRESETn VGND VGND VPWR VPWR _23091_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_243_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21853_ _21320_/X _21843_/X _21852_/X VGND VGND VPWR VPWR _21853_/X sky130_fd_sc_hd__a21bo_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20804_ _13145_/A VGND VGND VPWR VPWR _20804_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17450__A _14232_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24572_ _24537_/CLK _24572_/D HRESETn VGND VGND VPWR VPWR _24572_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16719__B1 _16364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21784_ _22387_/A _21782_/X _21783_/X VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__and3_4
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22068__A _21263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23522_/CLK _23523_/D VGND VGND VPWR VPWR _23523_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20735_ _24024_/Q VGND VGND VPWR VPWR _20735_/Y sky130_fd_sc_hd__inv_2
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16066__A _14420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _23454_/CLK _23454_/D VGND VGND VPWR VPWR _13414_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20666_ _14242_/Y _20646_/X _20637_/A _20665_/X VGND VGND VPWR VPWR _20667_/A sky130_fd_sc_hd__a211o_4
XFILLER_184_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22405_ _22402_/Y _22403_/X _22404_/X _13566_/A _22524_/B VGND VGND VPWR VPWR _22406_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19377__A _19085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20597_ _18887_/B _20596_/Y _20597_/C VGND VGND VPWR VPWR _20597_/X sky130_fd_sc_hd__and3_4
X_23385_ _23385_/CLK scl_oen_o_S5 VGND VGND VPWR VPWR _21005_/A sky130_fd_sc_hd__dfxtp_4
X_25124_ _25125_/CLK _14491_/X HRESETn VGND VGND VPWR VPWR _25124_/Q sky130_fd_sc_hd__dfrtp_4
X_22336_ _22335_/X VGND VGND VPWR VPWR _22336_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25055_ _24340_/CLK _14857_/X HRESETn VGND VGND VPWR VPWR _25055_/Q sky130_fd_sc_hd__dfrtp_4
X_22267_ _18300_/B _22267_/B VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__or2_4
XFILLER_133_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12020_ _25318_/Q _12019_/Y _25318_/Q _12019_/Y VGND VGND VPWR VPWR _12020_/X sky130_fd_sc_hd__a2bb2o_4
X_24006_ _23385_/CLK _24006_/D HRESETn VGND VGND VPWR VPWR _24006_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21218_ _21218_/A _21217_/X VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__or2_4
X_22198_ _21062_/A VGND VGND VPWR VPWR _22204_/A sky130_fd_sc_hd__buf_2
XFILLER_132_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21149_ _25493_/Q _13798_/B _25302_/Q _12068_/X VGND VGND VPWR VPWR _21149_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24573__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13971_ _13962_/X _13963_/X _13970_/X VGND VGND VPWR VPWR _13979_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__24502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15710_ _14386_/A _15709_/X VGND VGND VPWR VPWR _15710_/X sky130_fd_sc_hd__or2_4
XFILLER_74_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12922_ _12787_/Y _12927_/B _12875_/X VGND VGND VPWR VPWR _12922_/Y sky130_fd_sc_hd__a21oi_4
X_24908_ _24022_/CLK _24908_/D HRESETn VGND VGND VPWR VPWR _24908_/Q sky130_fd_sc_hd__dfrtp_4
X_16690_ _16689_/Y _16685_/X _16334_/X _16685_/X VGND VGND VPWR VPWR _16690_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16958__B1 _16166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15641_ _15626_/A VGND VGND VPWR VPWR _15641_/X sky130_fd_sc_hd__buf_2
XFILLER_234_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12853_ _12853_/A VGND VGND VPWR VPWR _12853_/Y sky130_fd_sc_hd__inv_2
X_24839_ _24889_/CLK _15830_/X HRESETn VGND VGND VPWR VPWR _24839_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_160_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23836_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15630__B1 _15629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11803_/X VGND VGND VPWR VPWR _11804_/X sky130_fd_sc_hd__buf_2
X_18360_ _18357_/Y _18361_/A _18359_/Y VGND VGND VPWR VPWR _18360_/Y sky130_fd_sc_hd__o21ai_4
XPHY_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15584_/A VGND VGND VPWR VPWR _15572_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_17_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _25520_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _22428_/A VGND VGND VPWR VPWR _12784_/Y sky130_fd_sc_hd__inv_2
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17242_/X _17301_/X _17311_/C VGND VGND VPWR VPWR _24369_/D sky130_fd_sc_hd__and3_4
XPHY_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14510_/B _14520_/X _14521_/Y _14522_/X VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__o22a_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _21135_/A _21135_/B VGND VGND VPWR VPWR _13786_/A sky130_fd_sc_hd__or2_4
X_18291_ _18282_/X _18285_/X _18290_/X VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__o21a_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17383__B1 _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17353_/A VGND VGND VPWR VPWR _17242_/X sky130_fd_sc_hd__buf_2
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14453_/Y _14451_/X _14400_/X _14451_/X VGND VGND VPWR VPWR _14454_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15394__C1 _15348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11666_/A VGND VGND VPWR VPWR _11666_/Y sky130_fd_sc_hd__inv_2
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13469_/A _13403_/X _13405_/C VGND VGND VPWR VPWR _13406_/C sky130_fd_sc_hd__and3_4
XANTENNA__21610__A _21564_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19124__B2 _19121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _17052_/Y _17074_/X _17076_/X _17170_/Y VGND VGND VPWR VPWR _17173_/X sky130_fd_sc_hd__a211o_4
X_14385_ _14385_/A _16378_/B _16378_/C _16378_/D VGND VGND VPWR VPWR _21348_/A sky130_fd_sc_hd__or4_4
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16124_ _16122_/Y _16123_/X _15963_/X _16123_/X VGND VGND VPWR VPWR _24707_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22425__B _22425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13336_ _13153_/X VGND VGND VPWR VPWR _13469_/A sky130_fd_sc_hd__buf_2
XFILLER_128_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16055_ _24732_/Q VGND VGND VPWR VPWR _16055_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13267_ _13267_/A VGND VGND VPWR VPWR _13267_/X sky130_fd_sc_hd__buf_2
XFILLER_142_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15006_ _15206_/A _16750_/A _15206_/A _16750_/A VGND VGND VPWR VPWR _15011_/A sky130_fd_sc_hd__a2bb2o_4
X_12218_ _12218_/A VGND VGND VPWR VPWR _12218_/Y sky130_fd_sc_hd__inv_2
X_13198_ _13198_/A _23924_/Q VGND VGND VPWR VPWR _13198_/X sky130_fd_sc_hd__or2_4
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19814_ _23620_/Q VGND VGND VPWR VPWR _19814_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12149_ _25479_/Q _12148_/Y _25479_/Q _12148_/Y VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19745_ _13258_/B VGND VGND VPWR VPWR _19745_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17254__B _17389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16957_ _16957_/A VGND VGND VPWR VPWR _16957_/X sky130_fd_sc_hd__buf_2
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22195__B1 _23980_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15908_ _15875_/Y VGND VGND VPWR VPWR _15908_/X sky130_fd_sc_hd__buf_2
X_19676_ _19675_/Y VGND VGND VPWR VPWR _19676_/X sky130_fd_sc_hd__buf_2
XFILLER_49_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16888_ _16887_/X VGND VGND VPWR VPWR _16888_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18627_ _16612_/A _24139_/Q _16612_/Y _18626_/Y VGND VGND VPWR VPWR _18627_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15839_ _12327_/Y _15835_/X _15767_/X _15838_/X VGND VGND VPWR VPWR _24833_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18558_ _18484_/B _18558_/B VGND VGND VPWR VPWR _18559_/A sky130_fd_sc_hd__or2_4
XFILLER_212_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17509_ _24306_/Q VGND VGND VPWR VPWR _17585_/D sky130_fd_sc_hd__inv_2
X_18489_ _18489_/A _18488_/X VGND VGND VPWR VPWR _18490_/B sky130_fd_sc_hd__nor2_4
XFILLER_33_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20520_ _20520_/A VGND VGND VPWR VPWR _20520_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15924__A1 _15694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20451_ _20451_/A VGND VGND VPWR VPWR _20451_/X sky130_fd_sc_hd__buf_2
XFILLER_165_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20382_ _20381_/Y _20377_/X _20034_/X _20364_/Y VGND VGND VPWR VPWR _23412_/D sky130_fd_sc_hd__a2bb2o_4
X_23170_ _24712_/Q _23296_/B VGND VGND VPWR VPWR _23170_/X sky130_fd_sc_hd__or2_4
XANTENNA__22670__A1 _21547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22670__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22121_ _22121_/A VGND VGND VPWR VPWR _22121_/X sky130_fd_sc_hd__buf_2
XANTENNA__11758__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18454__A1_N _23250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22052_ _22400_/A _22011_/Y _22018_/X _21520_/X _22051_/X VGND VGND VPWR VPWR _22053_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20433__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21003_ _20504_/A _23974_/Q _13982_/A VGND VGND VPWR VPWR _23974_/D sky130_fd_sc_hd__a21o_4
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19660__A _19652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19051__B1 _18999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22954_ _24572_/Q _22954_/B _22954_/C VGND VGND VPWR VPWR _22954_/X sky130_fd_sc_hd__and3_4
X_21905_ _21267_/A VGND VGND VPWR VPWR _22094_/A sky130_fd_sc_hd__buf_2
X_22885_ _22787_/X _22880_/Y _22881_/X _22884_/X VGND VGND VPWR VPWR _22885_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15612__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_233_0_HCLK clkbuf_7_116_0_HCLK/X VGND VGND VPWR VPWR _24012_/CLK sky130_fd_sc_hd__clkbuf_1
X_24624_ _24625_/CLK _16357_/X HRESETn VGND VGND VPWR VPWR _24624_/Q sky130_fd_sc_hd__dfrtp_4
X_21836_ _21654_/X _21835_/X _24229_/Q _21282_/X VGND VGND VPWR VPWR _21836_/X sky130_fd_sc_hd__o22a_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12977__A1 _12828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24555_ _24523_/CLK _16543_/X HRESETn VGND VGND VPWR VPWR _16542_/A sky130_fd_sc_hd__dfrtp_4
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21767_ _21648_/A _21767_/B VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__or2_4
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17365__B1 _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23506_ _24684_/CLK _23506_/D VGND VGND VPWR VPWR _20133_/A sky130_fd_sc_hd__dfxtp_4
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20718_ _22120_/A _20712_/Y _13137_/B VGND VGND VPWR VPWR _20718_/X sky130_fd_sc_hd__o21a_4
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24486_ _24674_/CLK _16724_/X HRESETn VGND VGND VPWR VPWR _16723_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21698_ _21693_/X _21696_/X _21697_/X VGND VGND VPWR VPWR _21698_/X sky130_fd_sc_hd__o21a_4
XFILLER_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ _23582_/CLK _20318_/X VGND VGND VPWR VPWR _23437_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20649_ _15470_/Y _20646_/X _20637_/X _20648_/X VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__a211o_4
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22110__B1 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14170_ _14155_/X _14169_/Y _14450_/A _14120_/X VGND VGND VPWR VPWR _14170_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23368_ VGND VGND VPWR VPWR _23368_/HI scl_o_S4 sky130_fd_sc_hd__conb_1
XANTENNA__18865__B1 _24579_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13121_ _13121_/A _13120_/Y _13121_/C VGND VGND VPWR VPWR _13121_/X sky130_fd_sc_hd__and3_4
X_25107_ _23970_/CLK _14542_/X HRESETn VGND VGND VPWR VPWR _25107_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22319_ _22171_/A _22319_/B _22318_/X VGND VGND VPWR VPWR _22319_/X sky130_fd_sc_hd__and3_4
X_23299_ _23299_/A _23289_/X _23299_/C _23298_/X VGND VGND VPWR VPWR _23299_/X sky130_fd_sc_hd__or4_4
XANTENNA__24754__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13052_ _12992_/Y _13052_/B VGND VGND VPWR VPWR _13061_/B sky130_fd_sc_hd__or2_4
X_25038_ _25043_/CLK _25038_/D HRESETn VGND VGND VPWR VPWR _14902_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12003_ _24107_/Q _12002_/X VGND VGND VPWR VPWR _12003_/X sky130_fd_sc_hd__and2_4
XANTENNA__20424__B1 _19817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17860_ _16920_/Y _16901_/Y _16937_/Y _17860_/D VGND VGND VPWR VPWR _17861_/D sky130_fd_sc_hd__or4_4
XFILLER_79_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16811_ _16810_/X VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__buf_2
XANTENNA__17074__B _17345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17791_ _16957_/X _17781_/X _17790_/X _17787_/B VGND VGND VPWR VPWR _17791_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21308__C _21308_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19530_ _22358_/B _19529_/X _11939_/X _19529_/X VGND VGND VPWR VPWR _23716_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13954_ _24980_/Q _13954_/B _13963_/B VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__or3_4
X_16742_ _16737_/Y VGND VGND VPWR VPWR _16762_/A sky130_fd_sc_hd__buf_2
XANTENNA__19042__B1 _18991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12905_ _12817_/A _12908_/B VGND VGND VPWR VPWR _12905_/X sky130_fd_sc_hd__or2_4
XFILLER_35_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16673_ _16685_/A VGND VGND VPWR VPWR _16673_/X sky130_fd_sc_hd__buf_2
X_19461_ _19460_/Y VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__buf_2
XFILLER_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21605__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13885_ _25252_/Q _13869_/X _21568_/A _13864_/X VGND VGND VPWR VPWR _13885_/X sky130_fd_sc_hd__o22a_4
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15603__B1 _11797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18412_ _24182_/Q VGND VGND VPWR VPWR _18471_/A sky130_fd_sc_hd__inv_2
XFILLER_222_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12836_ _12836_/A _12836_/B _12836_/C _12836_/D VGND VGND VPWR VPWR _12845_/C sky130_fd_sc_hd__or4_4
X_15624_ _15623_/Y _15621_/X _11834_/X _15621_/X VGND VGND VPWR VPWR _15624_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19392_ _19391_/X VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_62_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15555_ _16003_/A VGND VGND VPWR VPWR _22891_/B sky130_fd_sc_hd__buf_2
X_18343_ _18959_/A _18959_/B _18959_/A _18959_/B VGND VGND VPWR VPWR _24213_/D sky130_fd_sc_hd__a2bb2o_4
X_12767_ _22985_/A VGND VGND VPWR VPWR _12767_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14550_/A _14504_/X _20449_/A VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__o21a_4
XFILLER_230_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _11718_/A _11718_/B VGND VGND VPWR VPWR _13607_/A sky130_fd_sc_hd__or2_4
X_18274_ _18273_/Y _18270_/Y _16861_/X _18270_/Y VGND VGND VPWR VPWR _24228_/D sky130_fd_sc_hd__a2bb2o_4
X_15486_ _15486_/A VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__buf_2
X_12698_ _12680_/A _12685_/D _12697_/X VGND VGND VPWR VPWR _25421_/D sky130_fd_sc_hd__and3_4
XANTENNA__22436__A _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _25144_/Q VGND VGND VPWR VPWR _14437_/Y sky130_fd_sc_hd__inv_2
X_17225_ _17225_/A _17222_/X _17223_/X _17224_/X VGND VGND VPWR VPWR _17239_/B sky130_fd_sc_hd__or4_4
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16434__A _16434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22155__B _22155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17156_ _17064_/A VGND VGND VPWR VPWR _17160_/C sky130_fd_sc_hd__buf_2
X_14368_ _25165_/Q _14360_/X _25164_/Q _14365_/X VGND VGND VPWR VPWR _14368_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16107_ _16106_/Y _16104_/X _15950_/X _16104_/X VGND VGND VPWR VPWR _16107_/X sky130_fd_sc_hd__a2bb2o_4
X_13319_ _13356_/A _23921_/Q VGND VGND VPWR VPWR _13322_/B sky130_fd_sc_hd__or2_4
X_17087_ _17057_/A _17093_/A VGND VGND VPWR VPWR _17088_/B sky130_fd_sc_hd__or2_4
X_14299_ _25306_/Q _14299_/B _13532_/X VGND VGND VPWR VPWR _14303_/B sky130_fd_sc_hd__or3_4
XANTENNA__24495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16038_ _24739_/Q VGND VGND VPWR VPWR _16038_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15685__A3 _15656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22171__A _22171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_251_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13793__A _16464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22955__A2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17989_ _18227_/A _17980_/X _17988_/X VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__or3_4
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19728_ _11855_/A VGND VGND VPWR VPWR _19728_/X sky130_fd_sc_hd__buf_2
X_19659_ _19151_/A VGND VGND VPWR VPWR _19659_/X sky130_fd_sc_hd__buf_2
XANTENNA__13017__B _13017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16609__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15513__A _15503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22670_ _21547_/X _22669_/X _21550_/X _24873_/Q _21551_/X VGND VGND VPWR VPWR _22671_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_198_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12959__A1 _12855_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21621_ _21625_/A _21621_/B VGND VGND VPWR VPWR _21623_/B sky130_fd_sc_hd__or2_4
XANTENNA__18836__A2_N _18737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24340_ _24340_/CLK _17419_/X HRESETn VGND VGND VPWR VPWR _21008_/B sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_63_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24346_/CLK sky130_fd_sc_hd__clkbuf_1
X_21552_ _21547_/X _21549_/X _21550_/X _24723_/Q _21551_/X VGND VGND VPWR VPWR _21552_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20503_ _14286_/Y _20503_/B _20683_/A VGND VGND VPWR VPWR _20503_/X sky130_fd_sc_hd__and3_4
XFILLER_166_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24271_ _24272_/CLK _17875_/Y HRESETn VGND VGND VPWR VPWR _24271_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21483_ _21675_/A _19981_/Y VGND VGND VPWR VPWR _21483_/X sky130_fd_sc_hd__or2_4
XFILLER_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23222_ _15099_/A _23313_/B VGND VGND VPWR VPWR _23222_/X sky130_fd_sc_hd__or2_4
XANTENNA__24963__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20434_ _13385_/B VGND VGND VPWR VPWR _20434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13687__B _11890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23153_ _16750_/A _23016_/X _22903_/X VGND VGND VPWR VPWR _23153_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20365_ _20364_/Y VGND VGND VPWR VPWR _20365_/X sky130_fd_sc_hd__buf_2
XFILLER_228_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15125__A2 _15124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22104_ _14954_/A _22299_/B _21741_/A _22103_/X VGND VGND VPWR VPWR _22105_/C sky130_fd_sc_hd__a211o_4
X_20296_ _20295_/Y _20291_/X _20146_/A _20278_/Y VGND VGND VPWR VPWR _20296_/X sky130_fd_sc_hd__a2bb2o_4
X_23084_ _23020_/A _23074_/Y _23079_/X _23084_/D VGND VGND VPWR VPWR _23084_/X sky130_fd_sc_hd__or4_4
XFILLER_162_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22035_ _22028_/A _19950_/Y VGND VGND VPWR VPWR _22036_/C sky130_fd_sc_hd__or2_4
XFILLER_88_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17903__A _22003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23986_ _24003_/CLK _23984_/Q HRESETn VGND VGND VPWR VPWR _21013_/C sky130_fd_sc_hd__dfstp_4
XFILLER_17_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21425__A _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22937_ _24034_/Q _21296_/X _13658_/D _21320_/X VGND VGND VPWR VPWR _22938_/B sky130_fd_sc_hd__a22oi_4
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11951__A _19639_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _13670_/A _13670_/B VGND VGND VPWR VPWR _13671_/B sky130_fd_sc_hd__or2_4
XFILLER_232_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22868_ _22810_/A VGND VGND VPWR VPWR _22868_/X sky130_fd_sc_hd__buf_2
XFILLER_188_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ _12621_/A _12725_/A _12550_/Y _12729_/A VGND VGND VPWR VPWR _12621_/X sky130_fd_sc_hd__or4_4
X_24607_ _24602_/CLK _24607_/D HRESETn VGND VGND VPWR VPWR _15158_/A sky130_fd_sc_hd__dfrtp_4
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21819_ _21688_/A _21819_/B VGND VGND VPWR VPWR _21820_/C sky130_fd_sc_hd__or2_4
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22799_ _22799_/A _22799_/B _22510_/C VGND VGND VPWR VPWR _22799_/X sky130_fd_sc_hd__or3_4
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15340_ _15340_/A _15340_/B VGND VGND VPWR VPWR _15340_/X sky130_fd_sc_hd__or2_4
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12552_ _12550_/A _24867_/Q _12550_/Y _12551_/Y VGND VGND VPWR VPWR _12553_/D sky130_fd_sc_hd__o22a_4
X_24538_ _24989_/CLK _16587_/X HRESETn VGND VGND VPWR VPWR _24538_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21234__A1_N _15674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _15271_/A _15271_/B VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__or2_4
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _25449_/Q _12482_/Y VGND VGND VPWR VPWR _12485_/B sky130_fd_sc_hd__or2_4
X_24469_ _24430_/CLK _16765_/X HRESETn VGND VGND VPWR VPWR _16764_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _16040_/Y _24395_/Q _24742_/Q _17105_/A VGND VGND VPWR VPWR _17010_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _14221_/Y _14219_/X _13524_/X _14210_/A VGND VGND VPWR VPWR _25209_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14153_ _14153_/A VGND VGND VPWR VPWR _14153_/X sky130_fd_sc_hd__buf_2
X_13104_ _13104_/A _13104_/B _13103_/Y VGND VGND VPWR VPWR _25348_/D sky130_fd_sc_hd__and3_4
XANTENNA__23087__A _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14084_ _14013_/A _14074_/X _14066_/X _13998_/X _14075_/X VGND VGND VPWR VPWR _14084_/X
+ sky130_fd_sc_hd__a32o_4
X_18961_ _18974_/A VGND VGND VPWR VPWR _18961_/X sky130_fd_sc_hd__buf_2
X_13035_ _13049_/A _13031_/B _13034_/X VGND VGND VPWR VPWR _13036_/A sky130_fd_sc_hd__or3_4
X_17912_ _22009_/A _17911_/X _22009_/A _17911_/X VGND VGND VPWR VPWR _24262_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22937__A2 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18892_ _18891_/X VGND VGND VPWR VPWR _18893_/A sky130_fd_sc_hd__buf_2
XANTENNA__16077__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17843_ _17766_/A _17843_/B VGND VGND VPWR VPWR _17844_/C sky130_fd_sc_hd__or2_4
XFILLER_227_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15824__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16092__A3 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17774_ _17562_/X _17773_/X VGND VGND VPWR VPWR _17774_/X sky130_fd_sc_hd__or2_4
X_14986_ _25043_/Q VGND VGND VPWR VPWR _14986_/Y sky130_fd_sc_hd__inv_2
X_19513_ _19507_/Y VGND VGND VPWR VPWR _19513_/X sky130_fd_sc_hd__buf_2
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16725_ _24485_/Q VGND VGND VPWR VPWR _16725_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13937_ _13962_/C _13937_/B VGND VGND VPWR VPWR _13967_/C sky130_fd_sc_hd__or2_4
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24082__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22570__B1 _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11861__A _11861_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _19438_/A VGND VGND VPWR VPWR _19444_/X sky130_fd_sc_hd__buf_2
X_13868_ _25258_/Q _13866_/X _13861_/X _13867_/Y VGND VGND VPWR VPWR _13868_/X sky130_fd_sc_hd__a211o_4
X_16656_ _23303_/A _16655_/X _16294_/X _16655_/X VGND VGND VPWR VPWR _24514_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12819_ _12819_/A VGND VGND VPWR VPWR _12819_/Y sky130_fd_sc_hd__inv_2
X_15607_ _22805_/A _15602_/X _11805_/X _15602_/X VGND VGND VPWR VPWR _24914_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19375_ _19373_/Y _19369_/X _19308_/X _19374_/X VGND VGND VPWR VPWR _23770_/D sky130_fd_sc_hd__a2bb2o_4
X_13799_ _14415_/A _14484_/A VGND VGND VPWR VPWR _14264_/A sky130_fd_sc_hd__or2_4
X_16587_ _16586_/Y _16584_/X _16417_/X _16584_/X VGND VGND VPWR VPWR _16587_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18326_ _17710_/X _17713_/X _18325_/X VGND VGND VPWR VPWR _18326_/X sky130_fd_sc_hd__or3_4
X_15538_ _15544_/A VGND VGND VPWR VPWR _15538_/X sky130_fd_sc_hd__buf_2
XFILLER_231_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21070__A _15674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15469_ _14289_/X _24087_/Q _15450_/Y _13924_/C _15447_/A VGND VGND VPWR VPWR _15469_/X
+ sky130_fd_sc_hd__a32o_4
X_18257_ _18245_/X _18247_/X _13844_/A _24238_/Q _18248_/X VGND VGND VPWR VPWR _24238_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16164__A _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24676__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17208_ _24348_/Q VGND VGND VPWR VPWR _17389_/A sky130_fd_sc_hd__inv_2
XFILLER_175_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18188_ _13639_/X _18188_/B _18188_/C VGND VGND VPWR VPWR _18188_/X sky130_fd_sc_hd__and3_4
XANTENNA__24605__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17139_ _17139_/A _17139_/B VGND VGND VPWR VPWR _17139_/X sky130_fd_sc_hd__or2_4
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20150_ _20149_/X VGND VGND VPWR VPWR _20150_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20081_ _20093_/A VGND VGND VPWR VPWR _20081_/X sky130_fd_sc_hd__buf_2
XANTENNA__15508__A _15503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14412__A _14412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12341__A2 _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15815__B1 _11776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _24100_/CLK _23840_/D VGND VGND VPWR VPWR _18133_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_217_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23771_ _25077_/CLK _19372_/X VGND VGND VPWR VPWR _23771_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15830__A3 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20983_ _12158_/X _20982_/B VGND VGND VPWR VPWR _20983_/X sky130_fd_sc_hd__and2_4
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25510_ _23678_/CLK _11958_/X HRESETn VGND VGND VPWR VPWR _20007_/A sky130_fd_sc_hd__dfrtp_4
X_22722_ _24735_/Q _22425_/B _21121_/A _22721_/X VGND VGND VPWR VPWR _22722_/X sky130_fd_sc_hd__a211o_4
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23105__A2 _22444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25441_ _24283_/CLK _25441_/D HRESETn VGND VGND VPWR VPWR _12272_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22653_ _21295_/A _22651_/X _22121_/X _22652_/X VGND VGND VPWR VPWR _22654_/B sky130_fd_sc_hd__o22a_4
XFILLER_201_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21604_ _21604_/A _21603_/X VGND VGND VPWR VPWR _21604_/Y sky130_fd_sc_hd__nor2_4
X_25372_ _24824_/CLK _12990_/X HRESETn VGND VGND VPWR VPWR _21056_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_159_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22584_ _17861_/C _22443_/A _12288_/Y _21542_/A VGND VGND VPWR VPWR _22584_/X sky130_fd_sc_hd__o22a_4
X_24323_ _23534_/CLK _24323_/D HRESETn VGND VGND VPWR VPWR _17512_/A sky130_fd_sc_hd__dfrtp_4
X_21535_ _21535_/A VGND VGND VPWR VPWR _21714_/A sky130_fd_sc_hd__buf_2
XFILLER_223_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24254_ _25082_/CLK _17972_/X HRESETn VGND VGND VPWR VPWR _24254_/Q sky130_fd_sc_hd__dfrtp_4
X_21466_ _21473_/A VGND VGND VPWR VPWR _21466_/X sky130_fd_sc_hd__buf_2
XANTENNA__15897__A3 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_7_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__22804__A _22479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23205_ _23205_/A _23296_/B VGND VGND VPWR VPWR _23205_/X sky130_fd_sc_hd__or2_4
XFILLER_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20417_ _20408_/X _20404_/X _14248_/A _23397_/Q _20406_/X VGND VGND VPWR VPWR _20417_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_175_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24185_ _24189_/CLK _24185_/D HRESETn VGND VGND VPWR VPWR _24185_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21397_ _21246_/A VGND VGND VPWR VPWR _21412_/A sky130_fd_sc_hd__buf_2
XFILLER_162_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23136_ _22535_/B VGND VGND VPWR VPWR _23136_/X sky130_fd_sc_hd__buf_2
X_20348_ _20342_/X _19599_/D _11847_/A _22275_/A _20346_/X VGND VGND VPWR VPWR _23426_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20324__A _20323_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23067_ _17266_/A _22926_/X _12817_/A _22927_/X VGND VGND VPWR VPWR _23068_/B sky130_fd_sc_hd__a2bb2o_4
X_20279_ _20278_/Y VGND VGND VPWR VPWR _20279_/X sky130_fd_sc_hd__buf_2
XANTENNA__16059__B1 _15905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22018_ _24236_/Q _22595_/B _22062_/A _22017_/Y VGND VGND VPWR VPWR _22018_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14840_ _14840_/A VGND VGND VPWR VPWR _24005_/D sky130_fd_sc_hd__buf_2
XANTENNA__23354__B _23354_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14771_ _14783_/A _14785_/A _25065_/Q VGND VGND VPWR VPWR _14772_/C sky130_fd_sc_hd__and3_4
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _11710_/A _11710_/B _11889_/Y VGND VGND VPWR VPWR _11984_/C sky130_fd_sc_hd__o21a_4
X_23969_ _23970_/CLK _20618_/X HRESETn VGND VGND VPWR VPWR _23969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13722_ _13686_/Y VGND VGND VPWR VPWR _13722_/X sky130_fd_sc_hd__buf_2
X_16510_ _16510_/A VGND VGND VPWR VPWR _16510_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17490_ _24328_/Q VGND VGND VPWR VPWR _17490_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13653_ _13652_/X VGND VGND VPWR VPWR _14320_/A sky130_fd_sc_hd__buf_2
X_16441_ _15114_/Y _16438_/X _16066_/X _16438_/X VGND VGND VPWR VPWR _24592_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14992__A _14985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12604_ _25412_/Q VGND VGND VPWR VPWR _12729_/A sky130_fd_sc_hd__inv_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16372_ _24618_/Q VGND VGND VPWR VPWR _16372_/Y sky130_fd_sc_hd__inv_2
X_19160_ _19158_/Y _19159_/X _19091_/X _19159_/X VGND VGND VPWR VPWR _23847_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _25268_/Q VGND VGND VPWR VPWR _13584_/Y sky130_fd_sc_hd__inv_2
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15323_ _15355_/A _15323_/B _15323_/C VGND VGND VPWR VPWR _25012_/D sky130_fd_sc_hd__and3_4
X_18111_ _18036_/A _18111_/B VGND VGND VPWR VPWR _18112_/C sky130_fd_sc_hd__or2_4
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _12535_/A VGND VGND VPWR VPWR _12535_/Y sky130_fd_sc_hd__inv_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19091_ _19091_/A VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__buf_2
XFILLER_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15254_ _15253_/X VGND VGND VPWR VPWR _15254_/Y sky130_fd_sc_hd__inv_2
X_18042_ _18227_/A _18037_/X _18041_/X VGND VGND VPWR VPWR _18042_/X sky130_fd_sc_hd__or3_4
XFILLER_157_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12466_ _12247_/X _12440_/C _12411_/X _12462_/Y VGND VGND VPWR VPWR _12467_/A sky130_fd_sc_hd__a211o_4
XFILLER_157_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14205_ _13893_/X _24010_/Q VGND VGND VPWR VPWR _14205_/X sky130_fd_sc_hd__or2_4
X_15185_ _15184_/X VGND VGND VPWR VPWR _25043_/D sky130_fd_sc_hd__inv_2
XFILLER_172_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12397_ _12397_/A _12395_/A VGND VGND VPWR VPWR _12398_/C sky130_fd_sc_hd__or2_4
XFILLER_153_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14136_ _25229_/Q _14112_/X _14128_/C _14115_/B VGND VGND VPWR VPWR _14136_/X sky130_fd_sc_hd__o22a_4
XFILLER_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19993_ _19993_/A VGND VGND VPWR VPWR _19993_/X sky130_fd_sc_hd__buf_2
XFILLER_152_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14067_ _14064_/X VGND VGND VPWR VPWR _14068_/A sky130_fd_sc_hd__inv_2
X_18944_ _18944_/A VGND VGND VPWR VPWR _18944_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23032__B2 _21607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13018_ _13010_/X _13026_/D _13011_/A VGND VGND VPWR VPWR _13019_/C sky130_fd_sc_hd__o21a_4
X_18875_ _18875_/A VGND VGND VPWR VPWR _18876_/A sky130_fd_sc_hd__inv_2
XFILLER_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17826_ _16950_/Y _17820_/X _17790_/X _17823_/B VGND VGND VPWR VPWR _17827_/A sky130_fd_sc_hd__a211o_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23264__B _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21065__A _21064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ _17864_/A _16937_/Y _17757_/C _17757_/D VGND VGND VPWR VPWR _17761_/C sky130_fd_sc_hd__or4_4
X_14969_ _14969_/A VGND VGND VPWR VPWR _14969_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21346__A1 _24521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15063__A _15057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _16708_/A VGND VGND VPWR VPWR _16708_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17688_ _17522_/Y _17676_/B VGND VGND VPWR VPWR _17689_/C sky130_fd_sc_hd__nand2_4
XFILLER_207_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15025__B2 _24452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19427_ _19426_/Y _19422_/X _19402_/X _19422_/X VGND VGND VPWR VPWR _23752_/D sky130_fd_sc_hd__a2bb2o_4
X_16639_ _24516_/Q VGND VGND VPWR VPWR _16643_/A sky130_fd_sc_hd__inv_2
XFILLER_222_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24857__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22608__B _21450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12830__A2_N _24794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19358_ _19357_/Y _19353_/X _19246_/X _19353_/X VGND VGND VPWR VPWR _19358_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22846__A1 _16687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18309_ _18306_/X _18308_/X _18303_/X VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__o21a_4
X_19289_ _21904_/B _19286_/X _16885_/X _19286_/X VGND VGND VPWR VPWR _23801_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17722__B1 _21485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21320_ _21320_/A VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__buf_2
XANTENNA__13311__A _13228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22624__A _22624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_137_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _24252_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_191_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21251_ _14719_/Y VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__buf_2
XFILLER_116_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20202_ _23480_/Q VGND VGND VPWR VPWR _21783_/B sky130_fd_sc_hd__inv_2
XANTENNA__12562__A2 _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21182_ _21182_/A _20340_/Y VGND VGND VPWR VPWR _21183_/C sky130_fd_sc_hd__or2_4
XFILLER_116_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11766__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20133_ _20133_/A VGND VGND VPWR VPWR _20133_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19227__B1 _19226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20064_ _20064_/A VGND VGND VPWR VPWR _22086_/B sky130_fd_sc_hd__inv_2
X_24941_ _23408_/CLK _24941_/D HRESETn VGND VGND VPWR VPWR _11739_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24872_ _24872_/CLK _15760_/X HRESETn VGND VGND VPWR VPWR _24872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23823_ _23830_/CLK _23823_/D VGND VGND VPWR VPWR _18168_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15803__A3 _15562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _23754_/CLK _19423_/X VGND VGND VPWR VPWR _23754_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20964_/Y _20965_/Y _13676_/X VGND VGND VPWR VPWR _20966_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16213__B1 _11773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22705_/A VGND VGND VPWR VPWR _22737_/A sky130_fd_sc_hd__inv_2
XFILLER_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23190__A _23148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ _24206_/CLK _19621_/X VGND VGND VPWR VPWR _23685_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _24061_/Q _20896_/A VGND VGND VPWR VPWR _20897_/X sky130_fd_sc_hd__or2_4
XFILLER_198_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24598__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25424_ _25425_/CLK _25424_/D HRESETn VGND VGND VPWR VPWR _12563_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_186_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22636_ _22635_/X VGND VGND VPWR VPWR _22636_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25355_ _25358_/CLK _25355_/D HRESETn VGND VGND VPWR VPWR _12367_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22567_ _21060_/A _22566_/X VGND VGND VPWR VPWR _22567_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_33_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_66_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12320_ _12320_/A VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__inv_2
X_24306_ _24302_/CLK _24306_/D HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21513_/X _21517_/X _11692_/Y _21513_/X VGND VGND VPWR VPWR _21518_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_96_0_HCLK clkbuf_7_97_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_96_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25286_ _24233_/CLK _25286_/D HRESETn VGND VGND VPWR VPWR _13740_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22498_ _21129_/X VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__buf_2
XFILLER_155_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12251_ _12296_/A VGND VGND VPWR VPWR _12439_/A sky130_fd_sc_hd__buf_2
X_24237_ _24238_/CLK _24237_/D HRESETn VGND VGND VPWR VPWR _24237_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21449_ _21449_/A VGND VGND VPWR VPWR _23321_/A sky130_fd_sc_hd__buf_2
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16532__A _16532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12182_ _12181_/X VGND VGND VPWR VPWR _12182_/Y sky130_fd_sc_hd__inv_2
X_24168_ _24192_/CLK _24168_/D HRESETn VGND VGND VPWR VPWR _18434_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11761__B1 _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23119_ _23119_/A _23119_/B VGND VGND VPWR VPWR _23119_/X sky130_fd_sc_hd__or2_4
XANTENNA__25386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_16990_ _16990_/A VGND VGND VPWR VPWR _17072_/A sky130_fd_sc_hd__inv_2
X_24099_ _25106_/CLK _20478_/X HRESETn VGND VGND VPWR VPWR _24099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21555__A2_N _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15941_ _15940_/X VGND VGND VPWR VPWR _15941_/X sky130_fd_sc_hd__buf_2
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18459__A _18733_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18660_ _16576_/Y _24153_/Q _16606_/A _18794_/C VGND VGND VPWR VPWR _18660_/X sky130_fd_sc_hd__a2bb2o_4
X_15872_ _15871_/X VGND VGND VPWR VPWR _15872_/X sky130_fd_sc_hd__buf_2
XFILLER_209_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16452__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17611_ _17895_/B VGND VGND VPWR VPWR _17611_/X sky130_fd_sc_hd__buf_2
XFILLER_91_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14823_ _14823_/A _14823_/B _25052_/Q VGND VGND VPWR VPWR _14824_/B sky130_fd_sc_hd__or3_4
X_18591_ _18591_/A VGND VGND VPWR VPWR _18591_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17542_ _17542_/A _17542_/B _17540_/X _17542_/D VGND VGND VPWR VPWR _17542_/X sky130_fd_sc_hd__or4_4
X_11966_ _11656_/A VGND VGND VPWR VPWR _11967_/A sky130_fd_sc_hd__inv_2
X_14754_ _14753_/X VGND VGND VPWR VPWR _14755_/B sky130_fd_sc_hd__inv_2
XANTENNA__16204__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13705_ _13705_/A VGND VGND VPWR VPWR _13705_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14685_ _25068_/Q VGND VGND VPWR VPWR _14692_/A sky130_fd_sc_hd__buf_2
X_17473_ _18335_/A VGND VGND VPWR VPWR _18938_/B sky130_fd_sc_hd__buf_2
X_11897_ _11897_/A VGND VGND VPWR VPWR _11898_/A sky130_fd_sc_hd__inv_2
XANTENNA__24950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19212_ _19225_/A VGND VGND VPWR VPWR _19212_/X sky130_fd_sc_hd__buf_2
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22428__B _21091_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13636_ _13618_/X _14801_/A _13636_/C _13635_/X VGND VGND VPWR VPWR _13636_/X sky130_fd_sc_hd__or4_4
X_16424_ _16421_/Y _16423_/X _16334_/X _16423_/X VGND VGND VPWR VPWR _16424_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21332__B _21173_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19143_ _19143_/A _19143_/B _19346_/C VGND VGND VPWR VPWR _19143_/X sky130_fd_sc_hd__or3_4
X_13567_ _13566_/Y _14568_/A _13566_/Y _14568_/A VGND VGND VPWR VPWR _13567_/X sky130_fd_sc_hd__a2bb2o_4
X_16355_ _16354_/Y _16352_/X _16157_/X _16352_/X VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__a2bb2o_4
X_12518_ _12514_/A _12478_/B _12518_/C VGND VGND VPWR VPWR _25438_/D sky130_fd_sc_hd__and3_4
X_15306_ _15376_/A _15306_/B _15305_/X VGND VGND VPWR VPWR _15306_/X sky130_fd_sc_hd__or3_4
XFILLER_158_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16286_ _15678_/X _16288_/B _16090_/X _24649_/Q _16285_/X VGND VGND VPWR VPWR _16286_/X
+ sky130_fd_sc_hd__a32o_4
X_19074_ _23876_/Q VGND VGND VPWR VPWR _19074_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13498_ _13486_/A VGND VGND VPWR VPWR _13498_/X sky130_fd_sc_hd__buf_2
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22444__A _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18025_ _18168_/A _19214_/A VGND VGND VPWR VPWR _18026_/C sky130_fd_sc_hd__or2_4
X_12449_ _12208_/Y _12255_/Y _12197_/X _12449_/D VGND VGND VPWR VPWR _12449_/X sky130_fd_sc_hd__or4_4
X_15237_ _15252_/A _15232_/X _15236_/X VGND VGND VPWR VPWR _25030_/D sky130_fd_sc_hd__and3_4
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15191__B1 _15183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19457__B1 _19410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _15162_/Y VGND VGND VPWR VPWR _15310_/A sky130_fd_sc_hd__buf_2
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14119_ _14132_/B VGND VGND VPWR VPWR _14119_/X sky130_fd_sc_hd__buf_2
XFILLER_140_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16286__A3 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19753__A _11861_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15099_ _15099_/A VGND VGND VPWR VPWR _15099_/Y sky130_fd_sc_hd__inv_2
X_19976_ _19976_/A VGND VGND VPWR VPWR _19976_/Y sky130_fd_sc_hd__inv_2
X_18927_ _21773_/B _18922_/X _16890_/X _18922_/X VGND VGND VPWR VPWR _18927_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18858_ _16499_/Y _24150_/Q _16499_/Y _24150_/Q VGND VGND VPWR VPWR _18861_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16443__B1 _16070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17809_ _17753_/B _17803_/X _17790_/X _17805_/Y VGND VGND VPWR VPWR _17810_/A sky130_fd_sc_hd__a211o_4
XFILLER_54_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18789_ _18691_/B VGND VGND VPWR VPWR _18810_/A sky130_fd_sc_hd__buf_2
X_20820_ _20698_/X _20819_/Y _24926_/Q _20744_/A VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20751_ _20739_/X _20750_/Y _15616_/A _20744_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24691__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16617__A _16617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23470_ _25066_/CLK _23470_/D VGND VGND VPWR VPWR _23470_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20682_ _20686_/A _20682_/B VGND VGND VPWR VPWR _20682_/X sky130_fd_sc_hd__or2_4
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24620__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22421_ _22289_/X _22420_/X _21308_/C _16065_/A _21085_/X VGND VGND VPWR VPWR _22421_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_210_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16455__A2_N _16384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25140_ _25148_/CLK _25140_/D HRESETn VGND VGND VPWR VPWR _14450_/A sky130_fd_sc_hd__dfstp_4
X_22352_ _21945_/A _22350_/X _22351_/X VGND VGND VPWR VPWR _22352_/X sky130_fd_sc_hd__and3_4
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21303_ _21303_/A VGND VGND VPWR VPWR _21308_/C sky130_fd_sc_hd__buf_2
X_25071_ _25062_/CLK _25071_/D HRESETn VGND VGND VPWR VPWR _22055_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14459__A1_N _14186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22283_ _21588_/X VGND VGND VPWR VPWR _22283_/X sky130_fd_sc_hd__buf_2
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24022_ _24022_/CLK _24022_/D HRESETn VGND VGND VPWR VPWR _20725_/A sky130_fd_sc_hd__dfrtp_4
X_21234_ _15674_/A _21233_/X _13680_/Y _15674_/A VGND VGND VPWR VPWR _21234_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21165_ _21348_/B _21164_/X _17450_/B VGND VGND VPWR VPWR _21165_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17474__A2 _17461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20116_ _21791_/B _20109_/X _20115_/X _20109_/X VGND VGND VPWR VPWR _23512_/D sky130_fd_sc_hd__a2bb2o_4
X_21096_ _21592_/A VGND VGND VPWR VPWR _21096_/X sky130_fd_sc_hd__buf_2
XANTENNA__13496__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18279__A _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20047_ _20046_/Y _20044_/X _20000_/X _20044_/X VGND VGND VPWR VPWR _23537_/D sky130_fd_sc_hd__a2bb2o_4
X_24924_ _24923_/CLK _15582_/X HRESETn VGND VGND VPWR VPWR _15581_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24855_ _24878_/CLK _24855_/D HRESETn VGND VGND VPWR VPWR _24855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24779__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A VGND VGND VPWR VPWR _11820_/Y sky130_fd_sc_hd__inv_2
XPHY_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _25066_/CLK _19274_/X VGND VGND VPWR VPWR _23806_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24786_ _24787_/CLK _24786_/D HRESETn VGND VGND VPWR VPWR _24786_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _18277_/X _21985_/X _21989_/Y _22062_/A _21997_/X VGND VGND VPWR VPWR _21998_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24708__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22529__A _22529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11750_/X VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__buf_2
X_23737_ _23466_/CLK _19469_/X VGND VGND VPWR VPWR _18083_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_230_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _24073_/Q _20949_/B VGND VGND VPWR VPWR _20949_/X sky130_fd_sc_hd__or2_4
XPHY_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _25131_/Q VGND VGND VPWR VPWR _14470_/Y sky130_fd_sc_hd__inv_2
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _25300_/Q VGND VGND VPWR VPWR _11682_/Y sky130_fd_sc_hd__inv_2
X_23668_ _23916_/CLK _19678_/X VGND VGND VPWR VPWR _13158_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A _20095_/A VGND VGND VPWR VPWR _13422_/C sky130_fd_sc_hd__or2_4
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22619_ _21063_/A _22614_/X _21844_/X _22618_/Y VGND VGND VPWR VPWR _22620_/A sky130_fd_sc_hd__a211o_4
X_25407_ _25410_/CLK _12746_/X HRESETn VGND VGND VPWR VPWR _25407_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19687__B1 _19612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23494_/CLK _19875_/X VGND VGND VPWR VPWR _19873_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16140_ _16140_/A VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__inv_2
X_13352_ _13416_/A _13352_/B _13351_/X VGND VGND VPWR VPWR _13352_/X sky130_fd_sc_hd__or3_4
X_25338_ _25507_/CLK _25338_/D HRESETn VGND VGND VPWR VPWR _25338_/Q sky130_fd_sc_hd__dfrtp_4
X_12303_ _25371_/Q VGND VGND VPWR VPWR _13014_/A sky130_fd_sc_hd__inv_2
X_16071_ _16068_/Y _16069_/X _16070_/X _16069_/X VGND VGND VPWR VPWR _24727_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16595__A1_N _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13283_ _13322_/A _13283_/B _13282_/X VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__and3_4
X_25269_ _25281_/CLK _25269_/D HRESETn VGND VGND VPWR VPWR _13840_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17358__A _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15022_ _15022_/A VGND VGND VPWR VPWR _15022_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_120_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24042_/CLK sky130_fd_sc_hd__clkbuf_1
X_12234_ _25440_/Q _21544_/A _12232_/Y _12233_/Y VGND VGND VPWR VPWR _12235_/D sky130_fd_sc_hd__o22a_4
XFILLER_170_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_183_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _25148_/CLK sky130_fd_sc_hd__clkbuf_1
X_19830_ _19828_/Y _19829_/X _19734_/X _19829_/X VGND VGND VPWR VPWR _19830_/X sky130_fd_sc_hd__a2bb2o_4
X_12165_ _12101_/Y _12164_/X _12101_/Y _12164_/X VGND VGND VPWR VPWR _12166_/D sky130_fd_sc_hd__a2bb2o_4
X_19761_ _19761_/A VGND VGND VPWR VPWR _19761_/X sky130_fd_sc_hd__buf_2
X_12096_ _12094_/Y _12095_/X _11867_/X _12095_/X VGND VGND VPWR VPWR _12096_/X sky130_fd_sc_hd__a2bb2o_4
X_16973_ _16042_/Y _24394_/Q _16042_/Y _24394_/Q VGND VGND VPWR VPWR _16973_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13487__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18189__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18712_ _18720_/A _18717_/A _18711_/X VGND VGND VPWR VPWR _18712_/X sky130_fd_sc_hd__or3_4
X_15924_ _15694_/X _13597_/X _15701_/A _13551_/X VGND VGND VPWR VPWR _15924_/X sky130_fd_sc_hd__a211o_4
X_19692_ _19048_/A VGND VGND VPWR VPWR _19692_/X sky130_fd_sc_hd__buf_2
XFILLER_237_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12949__B _12609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18643_ _18643_/A _18623_/X _18632_/X _18642_/X VGND VGND VPWR VPWR _18643_/X sky130_fd_sc_hd__or4_4
X_15855_ _15664_/X _15774_/X _15851_/X _12613_/A _15854_/X VGND VGND VPWR VPWR _24823_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15325__B _15294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14806_ _14806_/A VGND VGND VPWR VPWR _14806_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17821__A _16950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18574_ _18479_/C _18573_/X _18494_/X VGND VGND VPWR VPWR _18574_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_92_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15786_ _15560_/X _15668_/B VGND VGND VPWR VPWR _15786_/X sky130_fd_sc_hd__or2_4
XFILLER_18_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _13068_/A _13063_/B _12998_/C VGND VGND VPWR VPWR _12998_/X sky130_fd_sc_hd__or3_4
XANTENNA__22439__A _22897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17525_ _17525_/A VGND VGND VPWR VPWR _17525_/Y sky130_fd_sc_hd__inv_2
X_14737_ _14736_/Y _14716_/Y _22055_/A _14715_/X VGND VGND VPWR VPWR _14749_/B sky130_fd_sc_hd__o22a_4
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11949_ _11947_/Y _11944_/X _11948_/X _11944_/X VGND VGND VPWR VPWR _11949_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23261__C _22954_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17456_ _17456_/A _11721_/Y _15791_/C _13476_/D VGND VGND VPWR VPWR _21178_/A sky130_fd_sc_hd__or4_4
XFILLER_220_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14668_ _14668_/A _14798_/A VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__or2_4
X_16407_ HWDATA[22] VGND VGND VPWR VPWR _16407_/X sky130_fd_sc_hd__buf_2
X_13619_ _13613_/B VGND VGND VPWR VPWR _18098_/A sky130_fd_sc_hd__buf_2
XFILLER_177_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19748__A _19742_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12214__A1 _25446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17387_ _17253_/Y _17390_/B _17280_/X VGND VGND VPWR VPWR _17387_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14599_ _14611_/A VGND VGND VPWR VPWR _14599_/X sky130_fd_sc_hd__buf_2
XFILLER_119_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19126_ _19134_/A VGND VGND VPWR VPWR _19126_/X sky130_fd_sc_hd__buf_2
XFILLER_158_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16338_ _16338_/A VGND VGND VPWR VPWR _16338_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17185__A2_N _17359_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20073__A2_N _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19057_ _19052_/Y _19056_/X _19032_/X _19056_/X VGND VGND VPWR VPWR _23884_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17268__A _17294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16269_ _16202_/A VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__buf_2
XANTENNA__16900__B2 _23332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18008_ _18008_/A VGND VGND VPWR VPWR _18126_/A sky130_fd_sc_hd__buf_2
XFILLER_160_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22902__A _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12205__A _21083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__A1 _14289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _21676_/B _19958_/X _19643_/X _19958_/X VGND VGND VPWR VPWR _23567_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22970_ _16733_/A _22967_/X _22969_/X VGND VGND VPWR VPWR _22970_/X sky130_fd_sc_hd__and3_4
XANTENNA__19602__B1 _19439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14420__A _14420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16416__B1 _16414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12859__B _12819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21921_ _21914_/A _21921_/B VGND VGND VPWR VPWR _21923_/B sky130_fd_sc_hd__or2_4
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24872__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24640_ _24641_/CLK _24640_/D HRESETn VGND VGND VPWR VPWR _16314_/A sky130_fd_sc_hd__dfrtp_4
X_21852_ _21124_/X _21846_/Y _21565_/A _21851_/X VGND VGND VPWR VPWR _21852_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24801__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20803_ _20788_/X _20802_/Y _15586_/A _20792_/X VGND VGND VPWR VPWR _24039_/D sky130_fd_sc_hd__a2bb2o_4
X_24571_ _24537_/CLK _24571_/D HRESETn VGND VGND VPWR VPWR _24571_/Q sky130_fd_sc_hd__dfrtp_4
X_21783_ _21783_/A _21783_/B VGND VGND VPWR VPWR _21783_/X sky130_fd_sc_hd__or2_4
XFILLER_224_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23522_ _23522_/CLK _20087_/X VGND VGND VPWR VPWR _13282_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ _20734_/A VGND VGND VPWR VPWR _20734_/Y sky130_fd_sc_hd__inv_2
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23913_/CLK _20275_/X VGND VGND VPWR VPWR _13446_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20665_ _17406_/B _20664_/Y _20669_/C VGND VGND VPWR VPWR _20665_/X sky130_fd_sc_hd__and3_4
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22404_ _22404_/A _21656_/X VGND VGND VPWR VPWR _22404_/X sky130_fd_sc_hd__or2_4
X_23384_ _23395_/CLK scl_oen_o_S4 VGND VGND VPWR VPWR _20987_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_136_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20596_ _23959_/Q _18886_/B VGND VGND VPWR VPWR _20596_/Y sky130_fd_sc_hd__nand2_4
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25123_ _25125_/CLK _14493_/X HRESETn VGND VGND VPWR VPWR _14492_/A sky130_fd_sc_hd__dfrtp_4
X_22335_ _14194_/Y _21861_/A _14263_/Y _14266_/A VGND VGND VPWR VPWR _22335_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25145__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16082__A _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25054_ _24340_/CLK _14860_/X HRESETn VGND VGND VPWR VPWR _25054_/Q sky130_fd_sc_hd__dfrtp_4
X_22266_ _22266_/A _22262_/X _22265_/X VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__or3_4
XANTENNA__22812__A _22811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24005_ _23980_/CLK _24005_/D HRESETn VGND VGND VPWR VPWR _24005_/Q sky130_fd_sc_hd__dfstp_4
X_21217_ _21217_/A _21351_/A VGND VGND VPWR VPWR _21217_/X sky130_fd_sc_hd__or2_4
X_22197_ _21350_/Y _22183_/X _22185_/X _22189_/Y _22196_/X VGND VGND VPWR VPWR _22205_/C
+ sky130_fd_sc_hd__a2111o_4
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22531__B _22531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21148_ _12108_/B _21146_/X _13504_/B _21147_/X VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__o22a_4
XFILLER_132_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13970_ _13969_/A _13968_/Y _13969_/Y _13967_/X VGND VGND VPWR VPWR _13970_/X sky130_fd_sc_hd__o22a_4
X_21079_ _21079_/A _21066_/X _21078_/X VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__and3_4
XFILLER_247_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20203__B2 _20198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12921_ _12773_/Y _12819_/Y _12921_/C _12921_/D VGND VGND VPWR VPWR _12927_/B sky130_fd_sc_hd__or4_4
X_24907_ _24022_/CLK _15624_/X HRESETn VGND VGND VPWR VPWR _15623_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20986__B _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18737__A _18737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ _24901_/Q VGND VGND VPWR VPWR _21757_/A sky130_fd_sc_hd__inv_2
XFILLER_246_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12852_ _25383_/Q VGND VGND VPWR VPWR _12855_/C sky130_fd_sc_hd__inv_2
X_24838_ _24883_/CLK _15831_/X HRESETn VGND VGND VPWR VPWR _24838_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23362__B _25175_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23153__B1 _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22259__A _21679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11803_ _11749_/X VGND VGND VPWR VPWR _11803_/X sky130_fd_sc_hd__buf_2
XANTENNA__19274__A2_N _19271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _25380_/Q VGND VGND VPWR VPWR _12783_/Y sky130_fd_sc_hd__inv_2
X_15571_ _15626_/A VGND VGND VPWR VPWR _15584_/A sky130_fd_sc_hd__buf_2
XPHY_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24757_/CLK _24769_/D HRESETn VGND VGND VPWR VPWR _22778_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17310_/A _17313_/B VGND VGND VPWR VPWR _17311_/C sky130_fd_sc_hd__or2_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _13822_/A _11734_/B VGND VGND VPWR VPWR _14417_/A sky130_fd_sc_hd__or2_4
X_14522_ _14510_/C VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__buf_2
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18290_ _18290_/A _20015_/B _18289_/X VGND VGND VPWR VPWR _18290_/X sky130_fd_sc_hd__or3_4
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16900__A2_N _23332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17240_/X VGND VGND VPWR VPWR _17353_/A sky130_fd_sc_hd__buf_2
XFILLER_230_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/A VGND VGND VPWR VPWR _13693_/A sky130_fd_sc_hd__inv_2
X_14453_ _25139_/Q VGND VGND VPWR VPWR _14453_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13372_/A _23615_/Q VGND VGND VPWR VPWR _13405_/C sky130_fd_sc_hd__or2_4
XFILLER_168_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19289__A2_N _19286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _13607_/A VGND VGND VPWR VPWR _14386_/A sky130_fd_sc_hd__buf_2
X_17172_ _17163_/X _17171_/X _17160_/C VGND VGND VPWR VPWR _17172_/X sky130_fd_sc_hd__and3_4
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13335_ _13254_/X _13333_/X _13334_/X VGND VGND VPWR VPWR _13335_/X sky130_fd_sc_hd__and3_4
X_16123_ _16103_/X VGND VGND VPWR VPWR _16123_/X sky130_fd_sc_hd__buf_2
XFILLER_155_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15697__A1 _15686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13266_ _13209_/X _13240_/X _13265_/X _25338_/Q _11974_/X VGND VGND VPWR VPWR _13266_/X
+ sky130_fd_sc_hd__o32a_4
X_16054_ _16053_/Y _16049_/X _11822_/X _16049_/X VGND VGND VPWR VPWR _24733_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15541__A2_N _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12217_ _25462_/Q _24777_/Q _12425_/A _12216_/Y VGND VGND VPWR VPWR _12221_/C sky130_fd_sc_hd__o22a_4
X_15005_ _14997_/X _14998_/X _15005_/C _15004_/X VGND VGND VPWR VPWR _15005_/X sky130_fd_sc_hd__or4_4
X_13197_ _13197_/A _13195_/X _13197_/C VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__and3_4
XFILLER_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19813_ _21247_/B _19806_/X _18934_/X _19788_/Y VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12148_ _12147_/X VGND VGND VPWR VPWR _12148_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21338__A _22171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11864__A _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19744_ _19740_/Y _19743_/X _19677_/X _19743_/X VGND VGND VPWR VPWR _19744_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12079_ _21580_/A VGND VGND VPWR VPWR _12080_/A sky130_fd_sc_hd__buf_2
X_16956_ _16100_/Y _24293_/Q _16100_/Y _24293_/Q VGND VGND VPWR VPWR _16956_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19857__A2_N _19851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15907_ _12794_/Y _15904_/X _15765_/X _15904_/X VGND VGND VPWR VPWR _15907_/X sky130_fd_sc_hd__a2bb2o_4
X_19675_ _19675_/A VGND VGND VPWR VPWR _19675_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16887_ _20119_/A VGND VGND VPWR VPWR _16887_/X sky130_fd_sc_hd__buf_2
X_18626_ _24139_/Q VGND VGND VPWR VPWR _18626_/Y sky130_fd_sc_hd__inv_2
X_15838_ _15806_/Y VGND VGND VPWR VPWR _15838_/X sky130_fd_sc_hd__buf_2
XFILLER_225_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18557_ _18488_/A _18557_/B VGND VGND VPWR VPWR _18558_/B sky130_fd_sc_hd__or2_4
XANTENNA__17270__B _17243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15769_ _12545_/Y _15763_/X _15767_/X _15768_/X VGND VGND VPWR VPWR _15769_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16167__A _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17508_ _11802_/Y _24312_/Q _11802_/Y _24312_/Q VGND VGND VPWR VPWR _17515_/A sky130_fd_sc_hd__a2bb2o_4
X_18488_ _18488_/A _18488_/B _18488_/C _18487_/X VGND VGND VPWR VPWR _18488_/X sky130_fd_sc_hd__or4_4
XFILLER_21_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14188__A1 _14186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21801__A _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _21733_/A _17434_/X _16796_/X _17434_/X VGND VGND VPWR VPWR _24334_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15385__B1 _15324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15924__A2 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20450_ _20448_/X _20451_/A VGND VGND VPWR VPWR _20469_/A sky130_fd_sc_hd__and2_4
XANTENNA__22655__C1 _22654_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19109_ _23864_/Q VGND VGND VPWR VPWR _21771_/B sky130_fd_sc_hd__inv_2
XFILLER_192_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20381_ _20381_/A VGND VGND VPWR VPWR _20381_/Y sky130_fd_sc_hd__inv_2
X_22120_ _22120_/A _21123_/A VGND VGND VPWR VPWR _22120_/X sky130_fd_sc_hd__or2_4
XFILLER_118_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22051_ _22274_/A _22030_/Y _22037_/Y _22044_/Y _22050_/Y VGND VGND VPWR VPWR _22051_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19823__B1 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21002_ _21002_/A _21002_/B VGND VGND VPWR VPWR _21002_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_23_0_HCLK clkbuf_8_23_0_HCLK/A VGND VGND VPWR VPWR _24715_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_229_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_86_0_HCLK clkbuf_8_86_0_HCLK/A VGND VGND VPWR VPWR _24849_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12769__A1_N _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14663__A2 _14650_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22953_ _16224_/A _22827_/B VGND VGND VPWR VPWR _22956_/B sky130_fd_sc_hd__or2_4
X_21904_ _22093_/A _21904_/B VGND VGND VPWR VPWR _21907_/B sky130_fd_sc_hd__or2_4
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22884_ _15800_/A _22883_/X _22503_/X _25543_/Q _22793_/X VGND VGND VPWR VPWR _22884_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21835_ _23423_/Q _20343_/X _23399_/Q _21972_/B VGND VGND VPWR VPWR _21835_/X sky130_fd_sc_hd__o22a_4
X_24623_ _24625_/CLK _24623_/D HRESETn VGND VGND VPWR VPWR _24623_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24554_ _24528_/CLK _16545_/X HRESETn VGND VGND VPWR VPWR _24554_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21766_ _21625_/A _21766_/B VGND VGND VPWR VPWR _21766_/X sky130_fd_sc_hd__or2_4
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17365__A1 _17359_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _13136_/A VGND VGND VPWR VPWR _22120_/A sky130_fd_sc_hd__inv_2
X_23505_ _23577_/CLK _23505_/D VGND VGND VPWR VPWR _23505_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24485_ _24485_/CLK _24485_/D HRESETn VGND VGND VPWR VPWR _24485_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21697_ _18301_/A VGND VGND VPWR VPWR _21697_/X sky130_fd_sc_hd__buf_2
XFILLER_168_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23436_ _23582_/CLK _20320_/X VGND VGND VPWR VPWR _20319_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20648_ _17402_/B _20648_/B _20628_/X VGND VGND VPWR VPWR _20648_/X sky130_fd_sc_hd__and3_4
XANTENNA__25159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22110__A1 _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23367_ VGND VGND VPWR VPWR _23367_/HI IRQ[31] sky130_fd_sc_hd__conb_1
XFILLER_165_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20579_ _20579_/A _18881_/X VGND VGND VPWR VPWR _20579_/Y sky130_fd_sc_hd__nand2_4
X_13120_ _12342_/Y _13115_/X VGND VGND VPWR VPWR _13120_/Y sky130_fd_sc_hd__nand2_4
X_22318_ _14931_/A _21341_/X _15676_/A _22317_/X VGND VGND VPWR VPWR _22318_/X sky130_fd_sc_hd__a211o_4
X_25106_ _25106_/CLK _14550_/X HRESETn VGND VGND VPWR VPWR scl_oen_o_S4 sky130_fd_sc_hd__dfstp_4
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23298_ _23123_/X _23295_/Y _23168_/X _23297_/X VGND VGND VPWR VPWR _23298_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13051_ _13051_/A VGND VGND VPWR VPWR _13069_/A sky130_fd_sc_hd__buf_2
X_25037_ _25043_/CLK _15210_/Y HRESETn VGND VGND VPWR VPWR _14927_/A sky130_fd_sc_hd__dfrtp_4
X_22249_ _22264_/A _19628_/Y VGND VGND VPWR VPWR _22250_/C sky130_fd_sc_hd__or2_4
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12002_ _24106_/Q _12001_/X VGND VGND VPWR VPWR _12002_/X sky130_fd_sc_hd__and2_4
XANTENNA__16628__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17355__B _17355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24794__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16810_ _16857_/A VGND VGND VPWR VPWR _16810_/X sky130_fd_sc_hd__buf_2
XANTENNA__15156__A _24605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19851__A _19838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17790_ _16963_/Y VGND VGND VPWR VPWR _17790_/X sky130_fd_sc_hd__buf_2
XANTENNA__24723__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12114__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16741_ _15026_/Y _16739_/X _15723_/X _16739_/X VGND VGND VPWR VPWR _16741_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23373__A _23360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13953_ _13952_/X VGND VGND VPWR VPWR _13953_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12904_ _12895_/X VGND VGND VPWR VPWR _12908_/B sky130_fd_sc_hd__inv_2
X_19460_ _19460_/A VGND VGND VPWR VPWR _19460_/Y sky130_fd_sc_hd__inv_2
X_16672_ _16653_/A VGND VGND VPWR VPWR _16685_/A sky130_fd_sc_hd__buf_2
X_13884_ _13880_/X _13883_/X _25194_/Q _13876_/X VGND VGND VPWR VPWR _13884_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17802__C _17562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18411_ _18411_/A _18406_/X _18411_/C _18411_/D VGND VGND VPWR VPWR _18430_/B sky130_fd_sc_hd__or4_4
XANTENNA__16800__B1 _16726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15623_ _15623_/A VGND VGND VPWR VPWR _15623_/Y sky130_fd_sc_hd__inv_2
X_12835_ _25395_/Q _12833_/Y _12834_/Y _24810_/Q VGND VGND VPWR VPWR _12836_/D sky130_fd_sc_hd__a2bb2o_4
X_19391_ _19391_/A VGND VGND VPWR VPWR _19391_/X sky130_fd_sc_hd__buf_2
XFILLER_222_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18342_ _18342_/A VGND VGND VPWR VPWR _18959_/B sky130_fd_sc_hd__buf_2
XFILLER_203_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15554_ _15553_/X VGND VGND VPWR VPWR _16003_/A sky130_fd_sc_hd__buf_2
X_12766_ _25383_/Q _12764_/Y _12765_/Y _23162_/A VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21152__A2 _24196_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _23941_/Q _23940_/Q VGND VGND VPWR VPWR _20449_/A sky130_fd_sc_hd__or2_4
XFILLER_15_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11717_ _13782_/A VGND VGND VPWR VPWR _11718_/B sky130_fd_sc_hd__inv_2
X_18273_ _18273_/A VGND VGND VPWR VPWR _18273_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15367__B1 _15324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _25421_/Q _12697_/B VGND VGND VPWR VPWR _12697_/X sky130_fd_sc_hd__or2_4
X_15485_ _15472_/A VGND VGND VPWR VPWR _15485_/X sky130_fd_sc_hd__buf_2
XFILLER_230_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16715__A _24489_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _16336_/Y _17340_/A _16336_/Y _17340_/A VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14436_ _14434_/Y _14435_/X _14404_/X _14435_/X VGND VGND VPWR VPWR _14436_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21340__B _22316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22101__B2 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _16969_/Y _17139_/X VGND VGND VPWR VPWR _17155_/Y sky130_fd_sc_hd__nand2_4
X_14367_ _14364_/X _14366_/Y _12072_/A _14364_/X VGND VGND VPWR VPWR _14367_/X sky130_fd_sc_hd__a2bb2o_4
X_16106_ _23237_/A VGND VGND VPWR VPWR _16106_/Y sky130_fd_sc_hd__inv_2
X_13318_ _13387_/A _13316_/X _13318_/C VGND VGND VPWR VPWR _13323_/B sky130_fd_sc_hd__and3_4
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14298_ _25184_/Q VGND VGND VPWR VPWR _14303_/A sky130_fd_sc_hd__inv_2
X_17086_ _17074_/A _17086_/B _17057_/B _17086_/D VGND VGND VPWR VPWR _17093_/A sky130_fd_sc_hd__or4_4
X_16037_ _16035_/Y _16031_/X _15967_/X _16036_/X VGND VGND VPWR VPWR _16037_/X sky130_fd_sc_hd__a2bb2o_4
X_13249_ _13249_/A _23795_/Q VGND VGND VPWR VPWR _13252_/B sky130_fd_sc_hd__or2_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16450__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16619__B1 _16534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13793__B _16464_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21068__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19761__A _19761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17988_ _17988_/A _17988_/B _17988_/C VGND VGND VPWR VPWR _17988_/X sky130_fd_sc_hd__and3_4
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19727_ _13333_/B VGND VGND VPWR VPWR _19727_/Y sky130_fd_sc_hd__inv_2
X_16939_ _16145_/Y _24275_/Q _16145_/Y _24275_/Q VGND VGND VPWR VPWR _16939_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13853__B1 _13809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19658_ _13292_/B VGND VGND VPWR VPWR _19658_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18609_ _16617_/A _18691_/B _16564_/Y _24158_/Q VGND VGND VPWR VPWR _18612_/C sky130_fd_sc_hd__a2bb2o_4
X_19589_ _23694_/Q VGND VGND VPWR VPWR _21505_/B sky130_fd_sc_hd__inv_2
XANTENNA__16807__A2_N _16806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21620_ _22226_/A VGND VGND VPWR VPWR _21625_/A sky130_fd_sc_hd__buf_2
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21531__A _21531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21551_ _21436_/X VGND VGND VPWR VPWR _21551_/X sky130_fd_sc_hd__buf_2
X_20502_ _20487_/A VGND VGND VPWR VPWR _20683_/A sky130_fd_sc_hd__buf_2
X_24270_ _24732_/CLK _17879_/X HRESETn VGND VGND VPWR VPWR _24270_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21482_ _21482_/A _21480_/X _21481_/X VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__and3_4
XANTENNA__25252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23221_ _23013_/A _23221_/B _23221_/C VGND VGND VPWR VPWR _23221_/X sky130_fd_sc_hd__and3_4
X_20433_ _20432_/Y _20430_/X _15777_/X _20430_/X VGND VGND VPWR VPWR _23390_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16858__B1 _16791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20654__A1 _14250_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23152_ _24610_/Q _23189_/B VGND VGND VPWR VPWR _23152_/X sky130_fd_sc_hd__or2_4
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20364_ _20364_/A VGND VGND VPWR VPWR _20364_/Y sky130_fd_sc_hd__inv_2
X_22103_ _24456_/Q _21091_/B _21344_/X VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__o21a_4
XFILLER_161_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14333__A1 _14338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083_ _22950_/A _23080_/X _23082_/X VGND VGND VPWR VPWR _23084_/D sky130_fd_sc_hd__and3_4
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20295_ _23445_/Q VGND VGND VPWR VPWR _20295_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22034_ _22034_/A _22034_/B VGND VGND VPWR VPWR _22036_/B sky130_fd_sc_hd__or2_4
XANTENNA__21603__B1 _22298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19272__B2 _19271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _24343_/CLK _23983_/Q HRESETn VGND VGND VPWR VPWR _23985_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__20610__A _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22936_ _23072_/A _22936_/B VGND VGND VPWR VPWR _22936_/Y sky130_fd_sc_hd__nor2_4
XFILLER_90_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22867_ _22866_/X VGND VGND VPWR VPWR _22867_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13224__A _13217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _12679_/A _12596_/Y _12620_/C VGND VGND VPWR VPWR _12628_/A sky130_fd_sc_hd__or3_4
X_24606_ _24602_/CLK _24606_/D HRESETn VGND VGND VPWR VPWR _15098_/A sky130_fd_sc_hd__dfrtp_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21818_ _21682_/A _21818_/B VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__or2_4
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22798_ _17262_/Y _22442_/A _25389_/Q _22306_/X VGND VGND VPWR VPWR _22799_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12551_ _24867_/Q VGND VGND VPWR VPWR _12551_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15349__B1 _15348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21441__A _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21749_ _22542_/A VGND VGND VPWR VPWR _21755_/A sky130_fd_sc_hd__buf_2
X_24537_ _24537_/CLK _16589_/X HRESETn VGND VGND VPWR VPWR _24537_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12481_/X VGND VGND VPWR VPWR _12482_/Y sky130_fd_sc_hd__inv_2
X_15270_ _15270_/A _15270_/B VGND VGND VPWR VPWR _15270_/X sky130_fd_sc_hd__or2_4
XANTENNA__22619__C1 _22618_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24468_ _24430_/CLK _24468_/D HRESETn VGND VGND VPWR VPWR _24468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _14221_/A VGND VGND VPWR VPWR _14221_/Y sky130_fd_sc_hd__inv_2
X_23419_ _23563_/CLK _20366_/X VGND VGND VPWR VPWR _20362_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24399_ _24406_/CLK _24399_/D HRESETn VGND VGND VPWR VPWR _24399_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22634__A2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14152_ _14119_/X _14151_/X _25145_/Q _14145_/X VGND VGND VPWR VPWR _14152_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_137_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25201__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _12326_/Y _13106_/B VGND VGND VPWR VPWR _13103_/Y sky130_fd_sc_hd__nand2_4
X_14083_ _20530_/A _14078_/X _14082_/X _14021_/B _14075_/X VGND VGND VPWR VPWR _14083_/X
+ sky130_fd_sc_hd__a32o_4
X_18960_ _18959_/X VGND VGND VPWR VPWR _18974_/A sky130_fd_sc_hd__inv_2
XANTENNA__15521__B1 HADDR[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23087__B _23087_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24904__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13034_ _13008_/X _13026_/D _13026_/A VGND VGND VPWR VPWR _13034_/X sky130_fd_sc_hd__o21a_4
X_17911_ _17913_/B _17908_/Y _17907_/X _17910_/X VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__o22a_4
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18891_ _18875_/A _18891_/B VGND VGND VPWR VPWR _18891_/X sky130_fd_sc_hd__or2_4
XFILLER_239_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17842_ _17764_/A _17842_/B VGND VGND VPWR VPWR _17844_/B sky130_fd_sc_hd__or2_4
XANTENNA__23347__B1 _22815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17773_ _16910_/Y _17793_/B VGND VGND VPWR VPWR _17773_/X sky130_fd_sc_hd__or2_4
XFILLER_208_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14985_ _14990_/A _24422_/Q _25014_/Q _14953_/Y VGND VGND VPWR VPWR _14985_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13835__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19512_ _23722_/Q VGND VGND VPWR VPWR _22022_/B sky130_fd_sc_hd__inv_2
XFILLER_235_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16724_ _16723_/Y _16721_/X _16451_/X _16721_/X VGND VGND VPWR VPWR _16724_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13936_ _13902_/A _13896_/A _13936_/C _13936_/D VGND VGND VPWR VPWR _13962_/C sky130_fd_sc_hd__or4_4
XFILLER_93_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19443_ _18044_/B VGND VGND VPWR VPWR _19443_/Y sky130_fd_sc_hd__inv_2
X_16655_ _16654_/X VGND VGND VPWR VPWR _16655_/X sky130_fd_sc_hd__buf_2
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867_ _13867_/A VGND VGND VPWR VPWR _13867_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15606_ _24914_/Q VGND VGND VPWR VPWR _22805_/A sky130_fd_sc_hd__inv_2
X_12818_ _12817_/Y _23054_/A _12817_/Y _23054_/A VGND VGND VPWR VPWR _12824_/B sky130_fd_sc_hd__a2bb2o_4
X_19374_ _19368_/Y VGND VGND VPWR VPWR _19374_/X sky130_fd_sc_hd__buf_2
XFILLER_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16586_ _24538_/Q VGND VGND VPWR VPWR _16586_/Y sky130_fd_sc_hd__inv_2
X_13798_ _21140_/A _13798_/B _17448_/A _17448_/B VGND VGND VPWR VPWR _14484_/A sky130_fd_sc_hd__or4_4
XFILLER_203_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18325_ _18325_/A _17743_/B _18322_/X _18324_/X VGND VGND VPWR VPWR _18325_/X sky130_fd_sc_hd__or4_4
XANTENNA__21351__A _21351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15537_ _21135_/A VGND VGND VPWR VPWR _15537_/Y sky130_fd_sc_hd__inv_2
X_12749_ _24785_/Q VGND VGND VPWR VPWR _12749_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18256_ _11695_/Y _18252_/X _16613_/X _18252_/X VGND VGND VPWR VPWR _24239_/D sky130_fd_sc_hd__a2bb2o_4
X_15468_ _13924_/C _20620_/A _15440_/X _13902_/A _15447_/A VGND VGND VPWR VPWR _15468_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13788__B _14228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17207_ _24626_/Q _24355_/Q _16351_/Y _17364_/A VGND VGND VPWR VPWR _17210_/C sky130_fd_sc_hd__o22a_4
XFILLER_163_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14419_ HWDATA[7] VGND VGND VPWR VPWR _14420_/A sky130_fd_sc_hd__buf_2
X_18187_ _18059_/A _18183_/X _18186_/X VGND VGND VPWR VPWR _18188_/C sky130_fd_sc_hd__or3_4
XANTENNA__19756__A _19742_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15760__B1 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _15399_/A _15398_/X VGND VGND VPWR VPWR _15399_/X sky130_fd_sc_hd__or2_4
XFILLER_156_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17138_ _17051_/Y _17138_/B VGND VGND VPWR VPWR _17139_/B sky130_fd_sc_hd__or2_4
XFILLER_190_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21833__B1 _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17276__A _17355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17069_ _17034_/X _17079_/A VGND VGND VPWR VPWR _17072_/B sky130_fd_sc_hd__or2_4
XFILLER_116_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24645__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20080_ _20079_/X VGND VGND VPWR VPWR _20093_/A sky130_fd_sc_hd__inv_2
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22910__A _22910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23770_ _25077_/CLK _23770_/D VGND VGND VPWR VPWR _23770_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20982_ _20982_/A _20982_/B VGND VGND VPWR VPWR _24117_/D sky130_fd_sc_hd__and2_4
XFILLER_226_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22721_ _16338_/A _22721_/B _21096_/X VGND VGND VPWR VPWR _22721_/X sky130_fd_sc_hd__and3_4
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22652_ _16699_/Y _22578_/B VGND VGND VPWR VPWR _22652_/X sky130_fd_sc_hd__and2_4
X_25440_ _24283_/CLK _25440_/D HRESETn VGND VGND VPWR VPWR _25440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14251__B1 _13819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21603_ _21606_/A _21600_/X _22298_/A _21602_/X VGND VGND VPWR VPWR _21603_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22583_ _21027_/X VGND VGND VPWR VPWR _22678_/B sky130_fd_sc_hd__buf_2
X_25371_ _25365_/CLK _13015_/X HRESETn VGND VGND VPWR VPWR _25371_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21534_ _21711_/A _21533_/X VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__and2_4
X_24322_ _23534_/CLK _17620_/Y HRESETn VGND VGND VPWR VPWR _24322_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24253_ _25082_/CLK _18032_/X HRESETn VGND VGND VPWR VPWR _24253_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21465_ _21210_/A VGND VGND VPWR VPWR _21473_/A sky130_fd_sc_hd__buf_2
X_23204_ _23203_/X VGND VGND VPWR VPWR _23204_/Y sky130_fd_sc_hd__inv_2
X_20416_ _20408_/X _20404_/X _20249_/X _23398_/Q _20406_/X VGND VGND VPWR VPWR _23398_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24184_ _24189_/CLK _24184_/D HRESETn VGND VGND VPWR VPWR _24184_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23188__A _22171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21396_ _21392_/X _21395_/X _21251_/X VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__o21a_4
XFILLER_119_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23135_ _23133_/X _23134_/X _22929_/X VGND VGND VPWR VPWR _23135_/X sky130_fd_sc_hd__or3_4
X_20347_ _20342_/X _19599_/D _13844_/A _21996_/A _20346_/X VGND VGND VPWR VPWR _23427_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16090__A _13818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23066_ _12424_/A _22998_/X _17751_/A _22924_/X VGND VGND VPWR VPWR _23066_/X sky130_fd_sc_hd__a2bb2o_4
X_20278_ _20278_/A VGND VGND VPWR VPWR _20278_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22017_ _22017_/A VGND VGND VPWR VPWR _22017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13219__A _13228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_56_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14770_ _14769_/X VGND VGND VPWR VPWR _14781_/A sky130_fd_sc_hd__inv_2
XFILLER_91_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11982_ _11661_/A _11981_/X _11979_/A _11890_/X VGND VGND VPWR VPWR _11985_/A sky130_fd_sc_hd__o22a_4
X_23968_ _23395_/CLK _20989_/X HRESETn VGND VGND VPWR VPWR _23968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13721_ _13698_/A _13698_/B VGND VGND VPWR VPWR _13721_/Y sky130_fd_sc_hd__nand2_4
XFILLER_216_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22919_ _22919_/A VGND VGND VPWR VPWR _22919_/Y sky130_fd_sc_hd__inv_2
X_23899_ _23880_/CLK _23899_/D VGND VGND VPWR VPWR _23899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16440_ _15108_/Y _16438_/X _16157_/X _16438_/X VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13652_ _13652_/A _14310_/A VGND VGND VPWR VPWR _13652_/X sky130_fd_sc_hd__or2_4
XANTENNA__25174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22304__A1 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12603_ _25434_/Q _12591_/Y _12590_/Y _24864_/Q VGND VGND VPWR VPWR _12603_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16371_ _16370_/Y _16365_/X _15995_/X _16365_/X VGND VGND VPWR VPWR _16371_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13583_ _25263_/Q _13582_/A _13581_/Y _13582_/Y VGND VGND VPWR VPWR _13587_/C sky130_fd_sc_hd__o22a_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22855__A2 _22851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12793__A _12793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _18072_/X _23768_/Q VGND VGND VPWR VPWR _18112_/B sky130_fd_sc_hd__or2_4
XFILLER_200_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15322_ _15322_/A _15319_/X VGND VGND VPWR VPWR _15323_/C sky130_fd_sc_hd__or2_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12534_ _12622_/A _12532_/Y _12630_/A _24886_/Q VGND VGND VPWR VPWR _12534_/X sky130_fd_sc_hd__a2bb2o_4
X_19090_ _19090_/A VGND VGND VPWR VPWR _19090_/X sky130_fd_sc_hd__buf_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18041_ _17988_/A _18039_/X _18040_/X VGND VGND VPWR VPWR _18041_/X sky130_fd_sc_hd__and3_4
X_15253_ _15248_/A _15247_/X _15208_/X _15249_/Y VGND VGND VPWR VPWR _15253_/X sky130_fd_sc_hd__a211o_4
X_12465_ _12458_/A _12463_/X _12465_/C VGND VGND VPWR VPWR _25453_/D sky130_fd_sc_hd__and3_4
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15742__B1 _11787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14204_ _14204_/A _14203_/X VGND VGND VPWR VPWR _14207_/B sky130_fd_sc_hd__or2_4
X_12396_ _12188_/A _12395_/Y VGND VGND VPWR VPWR _12398_/B sky130_fd_sc_hd__or2_4
X_15184_ _14986_/Y _15182_/X _15183_/X _15176_/Y VGND VGND VPWR VPWR _15184_/X sky130_fd_sc_hd__a211o_4
XFILLER_172_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14135_ _14117_/X VGND VGND VPWR VPWR _14141_/A sky130_fd_sc_hd__buf_2
X_19992_ _23555_/Q VGND VGND VPWR VPWR _22256_/B sky130_fd_sc_hd__inv_2
X_14066_ _14066_/A VGND VGND VPWR VPWR _14066_/X sky130_fd_sc_hd__buf_2
X_18943_ _18942_/Y _18940_/X _17430_/X _18940_/X VGND VGND VPWR VPWR _23923_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23032__A2 _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22730__A _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14232__B _14232_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21723__A2_N _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13017_ _13021_/C _13017_/B VGND VGND VPWR VPWR _13026_/D sky130_fd_sc_hd__and2_4
X_18874_ _18873_/X VGND VGND VPWR VPWR _18874_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21594__A2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18995__B1 _18975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17825_ _17852_/A _17823_/X _17825_/C VGND VGND VPWR VPWR _17825_/X sky130_fd_sc_hd__and3_4
XFILLER_227_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12968__A _12952_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17756_ _21066_/A VGND VGND VPWR VPWR _17757_/D sky130_fd_sc_hd__inv_2
XFILLER_208_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14968_ _15232_/A _14950_/A _14912_/X _14913_/Y VGND VGND VPWR VPWR _14972_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21346__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16707_ _16706_/Y _16704_/X _16609_/X _16704_/X VGND VGND VPWR VPWR _16707_/X sky130_fd_sc_hd__a2bb2o_4
X_13919_ _13937_/B VGND VGND VPWR VPWR _13927_/C sky130_fd_sc_hd__inv_2
XFILLER_235_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17687_ _17687_/A _17684_/B _17687_/C VGND VGND VPWR VPWR _17687_/X sky130_fd_sc_hd__and3_4
XFILLER_208_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14899_ _24425_/Q VGND VGND VPWR VPWR _14899_/Y sky130_fd_sc_hd__inv_2
X_19426_ _18117_/B VGND VGND VPWR VPWR _19426_/Y sky130_fd_sc_hd__inv_2
X_16638_ _24517_/Q VGND VGND VPWR VPWR _16640_/A sky130_fd_sc_hd__inv_2
XFILLER_23_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17970__A1 _15686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21081__A _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _18128_/B VGND VGND VPWR VPWR _19357_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16569_ _24545_/Q VGND VGND VPWR VPWR _16569_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15981__B1 _22644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18308_ _18310_/B _18301_/B VGND VGND VPWR VPWR _18308_/X sky130_fd_sc_hd__and2_4
XANTENNA__12795__B1 _12855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19288_ _23801_/Q VGND VGND VPWR VPWR _21904_/B sky130_fd_sc_hd__inv_2
XFILLER_175_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24897__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18239_ _17458_/C VGND VGND VPWR VPWR _20405_/A sky130_fd_sc_hd__buf_2
XANTENNA__24826__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21250_ _21638_/A _21250_/B _21250_/C VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__and3_4
XFILLER_117_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20201_ _20200_/Y _20198_/X _20112_/X _20198_/X VGND VGND VPWR VPWR _23481_/D sky130_fd_sc_hd__a2bb2o_4
X_21181_ _24217_/Q _21181_/B VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__or2_4
XANTENNA__14423__A _14423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20132_ _20131_/Y _20129_/X _20105_/X _20129_/X VGND VGND VPWR VPWR _20132_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20063_ _20062_/Y _20060_/X _19793_/X _20060_/X VGND VGND VPWR VPWR _20063_/X sky130_fd_sc_hd__a2bb2o_4
X_24940_ _23716_/CLK _15531_/X HRESETn VGND VGND VPWR VPWR _11739_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_246_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24871_ _24872_/CLK _24871_/D HRESETn VGND VGND VPWR VPWR _24871_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12384__A2_N _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23822_ _23830_/CLK _19229_/X VGND VGND VPWR VPWR _23822_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21337__A2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20965_ _20961_/X VGND VGND VPWR VPWR _20965_/Y sky130_fd_sc_hd__inv_2
X_23753_ _23754_/CLK _19425_/X VGND VGND VPWR VPWR _18080_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_213_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18565__A _18515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _22479_/A _22700_/X _23008_/A _22703_/X VGND VGND VPWR VPWR _22705_/A sky130_fd_sc_hd__o22a_4
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20896_/A VGND VGND VPWR VPWR _20896_/Y sky130_fd_sc_hd__inv_2
X_23684_ _23684_/CLK _23684_/D VGND VGND VPWR VPWR _23684_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14224__B1 _13819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15567__A3 _15562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15421__C1 _15348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22087__A _22387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25423_ _25425_/CLK _12693_/X HRESETn VGND VGND VPWR VPWR _12583_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22635_ _22528_/X _22632_/X _22431_/X _22634_/X VGND VGND VPWR VPWR _22635_/X sky130_fd_sc_hd__o22a_4
XFILLER_241_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22566_ _22563_/X _22564_/X _22145_/C _24870_/Q _22565_/X VGND VGND VPWR VPWR _22566_/X
+ sky130_fd_sc_hd__a32o_4
X_25354_ _25358_/CLK _13078_/Y HRESETn VGND VGND VPWR VPWR _12358_/A sky130_fd_sc_hd__dfrtp_4
X_21517_ _21514_/X _21383_/A _21517_/C VGND VGND VPWR VPWR _21517_/X sky130_fd_sc_hd__and3_4
X_24305_ _24302_/CLK _17685_/X HRESETn VGND VGND VPWR VPWR _24305_/Q sky130_fd_sc_hd__dfrtp_4
X_22497_ _21314_/A VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__buf_2
X_25285_ _23690_/CLK _13765_/Y HRESETn VGND VGND VPWR VPWR _25285_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24567__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12250_ _12250_/A VGND VGND VPWR VPWR _12296_/A sky130_fd_sc_hd__inv_2
X_21448_ _21081_/A VGND VGND VPWR VPWR _21449_/A sky130_fd_sc_hd__buf_2
X_24236_ _24238_/CLK _24236_/D HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23262__A2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11957__A _19639_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _13484_/C _12081_/B _13542_/C _12109_/A VGND VGND VPWR VPWR _12181_/X sky130_fd_sc_hd__or4_4
X_24167_ _24192_/CLK _18591_/Y HRESETn VGND VGND VPWR VPWR _24167_/Q sky130_fd_sc_hd__dfrtp_4
X_21379_ _21350_/Y _21361_/X _21367_/Y _21378_/Y VGND VGND VPWR VPWR _21425_/C sky130_fd_sc_hd__a211o_4
XFILLER_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23118_ _21535_/A VGND VGND VPWR VPWR _23118_/X sky130_fd_sc_hd__buf_2
XFILLER_162_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24098_ _25106_/CLK _20469_/X HRESETn VGND VGND VPWR VPWR _24098_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15940_ _15939_/X VGND VGND VPWR VPWR _15940_/X sky130_fd_sc_hd__buf_2
X_23049_ _23049_/A _23158_/B VGND VGND VPWR VPWR _23049_/X sky130_fd_sc_hd__or2_4
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22773__A1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15871_ _15896_/A VGND VGND VPWR VPWR _15871_/X sky130_fd_sc_hd__buf_2
XFILLER_49_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23084__C _23079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17610_ _17610_/A _17610_/B _17569_/B _17610_/D VGND VGND VPWR VPWR _17610_/X sky130_fd_sc_hd__or4_4
X_14822_ _24006_/Q _14822_/B _14822_/C VGND VGND VPWR VPWR _14823_/B sky130_fd_sc_hd__or3_4
XANTENNA__16452__B2 _16446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18590_ _18480_/Y _18566_/X _18588_/B _18505_/X VGND VGND VPWR VPWR _18591_/A sky130_fd_sc_hd__a211o_4
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17541_ _11811_/Y _24310_/Q _11811_/Y _24310_/Q VGND VGND VPWR VPWR _17542_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23381__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14753_ _14730_/C _14712_/A _14713_/Y VGND VGND VPWR VPWR _14753_/X sky130_fd_sc_hd__o21a_4
X_11965_ _11963_/Y _11956_/X _11964_/X _11934_/X VGND VGND VPWR VPWR _25508_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13704_ _24225_/Q _13703_/X VGND VGND VPWR VPWR _13705_/A sky130_fd_sc_hd__and2_4
XFILLER_189_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_143_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _23644_/CLK sky130_fd_sc_hd__clkbuf_1
X_17472_ _18332_/A VGND VGND VPWR VPWR _18335_/A sky130_fd_sc_hd__inv_2
XFILLER_72_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14684_ _14684_/A _11718_/B _13606_/X _13607_/B VGND VGND VPWR VPWR _14713_/A sky130_fd_sc_hd__or4_4
XANTENNA__14215__B1 _13849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11896_ _11933_/A _17711_/D _11881_/X _11891_/X _11895_/Y VGND VGND VPWR VPWR _11898_/B
+ sky130_fd_sc_hd__a2111o_4
XFILLER_220_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19211_ _19210_/X VGND VGND VPWR VPWR _19225_/A sky130_fd_sc_hd__buf_2
X_16423_ _16442_/A VGND VGND VPWR VPWR _16423_/X sky130_fd_sc_hd__buf_2
XFILLER_71_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13635_ _13634_/X _13635_/B VGND VGND VPWR VPWR _13635_/X sky130_fd_sc_hd__and2_4
XFILLER_204_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19142_ _13626_/A _19142_/B _14668_/A VGND VGND VPWR VPWR _19346_/C sky130_fd_sc_hd__or3_4
X_16354_ _24625_/Q VGND VGND VPWR VPWR _16354_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13566_ _13566_/A VGND VGND VPWR VPWR _13566_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22725__A _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ _15305_/A _15380_/A _15370_/A _15139_/Y VGND VGND VPWR VPWR _15305_/X sky130_fd_sc_hd__or4_4
X_12517_ _21083_/A _13049_/A VGND VGND VPWR VPWR _12518_/C sky130_fd_sc_hd__or2_4
X_19073_ _19072_/Y _19068_/X _18999_/X _19061_/A VGND VGND VPWR VPWR _23877_/D sky130_fd_sc_hd__a2bb2o_4
X_16285_ _16284_/X _16001_/X VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__or2_4
X_13497_ _13497_/A VGND VGND VPWR VPWR _13497_/Y sky130_fd_sc_hd__inv_2
X_18024_ _18013_/A VGND VGND VPWR VPWR _18168_/A sky130_fd_sc_hd__buf_2
X_15236_ _25030_/Q _15235_/Y VGND VGND VPWR VPWR _15236_/X sky130_fd_sc_hd__or2_4
X_12448_ _12447_/X VGND VGND VPWR VPWR _25458_/D sky130_fd_sc_hd__inv_2
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ _24987_/Q VGND VGND VPWR VPWR _15415_/A sky130_fd_sc_hd__inv_2
XANTENNA__22461__B1 _14925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12379_ _12370_/A _12377_/Y _13054_/A _24845_/Q VGND VGND VPWR VPWR _12380_/D sky130_fd_sc_hd__a2bb2o_4
X_14118_ _14117_/X VGND VGND VPWR VPWR _14132_/B sky130_fd_sc_hd__inv_2
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15098_ _15098_/A VGND VGND VPWR VPWR _15098_/Y sky130_fd_sc_hd__inv_2
X_19975_ _19974_/Y _19972_/X _19636_/X _19972_/X VGND VGND VPWR VPWR _19975_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22460__A _23087_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14049_ _13998_/X _14048_/Y _14021_/D _14022_/A VGND VGND VPWR VPWR _14050_/A sky130_fd_sc_hd__or4_4
X_18926_ _18926_/A VGND VGND VPWR VPWR _21773_/B sky130_fd_sc_hd__inv_2
XANTENNA__23275__B _22968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22764__B2 _22940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18857_ _16490_/Y _18744_/A _16490_/Y _18744_/A VGND VGND VPWR VPWR _18861_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17808_ _17748_/X _17806_/X _17807_/X VGND VGND VPWR VPWR _24288_/D sky130_fd_sc_hd__and3_4
X_18788_ _18626_/Y VGND VGND VPWR VPWR _18799_/B sky130_fd_sc_hd__buf_2
XANTENNA__25096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14454__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21226__D _21225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17739_ _24224_/Q VGND VGND VPWR VPWR _17740_/A sky130_fd_sc_hd__inv_2
XANTENNA__25025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19393__B1 _19326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20750_ _13141_/A _13140_/X _20749_/Y VGND VGND VPWR VPWR _20750_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_211_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15802__A _15802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19409_ _18207_/B VGND VGND VPWR VPWR _19409_/Y sky130_fd_sc_hd__inv_2
X_20681_ _20681_/A _14291_/X VGND VGND VPWR VPWR _20683_/B sky130_fd_sc_hd__or2_4
XANTENNA__15954__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14418__A _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22420_ _24624_/Q _22284_/X VGND VGND VPWR VPWR _22420_/X sky130_fd_sc_hd__or2_4
XANTENNA__13322__A _13322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22351_ _21938_/A _22351_/B VGND VGND VPWR VPWR _22351_/X sky130_fd_sc_hd__or2_4
XFILLER_164_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24660__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21302_ _22202_/C VGND VGND VPWR VPWR _21303_/A sky130_fd_sc_hd__buf_2
X_25070_ _25062_/CLK _25070_/D HRESETn VGND VGND VPWR VPWR _22056_/A sky130_fd_sc_hd__dfrtp_4
X_22282_ _21293_/X VGND VGND VPWR VPWR _22294_/A sky130_fd_sc_hd__buf_2
XFILLER_145_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15721__A3 _15562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24021_ _24022_/CLK _24021_/D HRESETn VGND VGND VPWR VPWR _24021_/Q sky130_fd_sc_hd__dfrtp_4
X_21233_ _21026_/B _16280_/A _15663_/X _20830_/A _15667_/A VGND VGND VPWR VPWR _21233_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21164_ _21157_/X _21164_/B _21162_/X _21164_/D VGND VGND VPWR VPWR _21164_/X sky130_fd_sc_hd__and4_4
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16131__B1 _15970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20115_ _20115_/A VGND VGND VPWR VPWR _20115_/X sky130_fd_sc_hd__buf_2
XFILLER_59_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21095_ _21048_/X _21094_/Y _24785_/Q _21048_/X VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__a2bb2o_4
X_20046_ _23537_/Q VGND VGND VPWR VPWR _20046_/Y sky130_fd_sc_hd__inv_2
X_24923_ _24923_/CLK _15585_/X HRESETn VGND VGND VPWR VPWR _15583_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24854_ _25425_/CLK _24854_/D HRESETn VGND VGND VPWR VPWR _24854_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25105__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23445_/CLK _23805_/D VGND VGND VPWR VPWR _19275_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21714__A _21714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24785_ _24787_/CLK _15937_/X HRESETn VGND VGND VPWR VPWR _24785_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _21993_/Y _21994_/X _21995_/X _21996_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__a211o_4
XPHY_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11749_/X VGND VGND VPWR VPWR _11750_/X sky130_fd_sc_hd__buf_2
X_23736_ _23466_/CLK _19471_/X VGND VGND VPWR VPWR _19470_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16198__B1 _11752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20949_/B VGND VGND VPWR VPWR _20948_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_216_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24562_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18852__A1_N _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _25301_/Q _22745_/A _11666_/A _22595_/A VGND VGND VPWR VPWR _11684_/C sky130_fd_sc_hd__a2bb2o_4
X_23667_ _23642_/CLK _23667_/D VGND VGND VPWR VPWR _19679_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _13670_/B VGND VGND VPWR VPWR _20879_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21740__A1_N _16271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24748__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13420_/A _23918_/Q VGND VGND VPWR VPWR _13422_/B sky130_fd_sc_hd__or2_4
X_25406_ _25410_/CLK _12748_/Y HRESETn VGND VGND VPWR VPWR _12538_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _22768_/A _22618_/B VGND VGND VPWR VPWR _22618_/Y sky130_fd_sc_hd__nor2_4
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23598_ _23597_/CLK _23598_/D VGND VGND VPWR VPWR _19876_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13351_ _13310_/X _13349_/X _13351_/C VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__and3_4
X_25337_ _25488_/CLK _13268_/X HRESETn VGND VGND VPWR VPWR _25337_/Q sky130_fd_sc_hd__dfrtp_4
X_22549_ _13589_/Y _22549_/B VGND VGND VPWR VPWR _22549_/X sky130_fd_sc_hd__and2_4
XFILLER_10_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11982__A1 _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12302_ _13002_/C _24836_/Q _13002_/C _24836_/Q VGND VGND VPWR VPWR _12310_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11982__B2 _11890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16070_ _14423_/A VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__buf_2
X_13282_ _13282_/A _13282_/B VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__or2_4
X_25268_ _25281_/CLK _25268_/D HRESETn VGND VGND VPWR VPWR _25268_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17358__B _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15021_ _15013_/X _15021_/B _15021_/C _15021_/D VGND VGND VPWR VPWR _15021_/X sky130_fd_sc_hd__or4_4
X_12233_ _21544_/A VGND VGND VPWR VPWR _12233_/Y sky130_fd_sc_hd__inv_2
X_24219_ _24217_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
X_25199_ _23998_/CLK _14251_/X HRESETn VGND VGND VPWR VPWR _25199_/Q sky130_fd_sc_hd__dfstp_4
X_12164_ _12160_/A _12157_/A _12162_/Y VGND VGND VPWR VPWR _12164_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23376__A _21002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12095_ _12083_/A VGND VGND VPWR VPWR _12095_/X sky130_fd_sc_hd__buf_2
X_16972_ _16967_/X _16972_/B _16970_/X _16972_/D VGND VGND VPWR VPWR _16972_/X sky130_fd_sc_hd__or4_4
X_19760_ _13465_/B VGND VGND VPWR VPWR _19760_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15923_ _13547_/A _15923_/B VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__and2_4
X_18711_ _18711_/A _18710_/X VGND VGND VPWR VPWR _18711_/X sky130_fd_sc_hd__or2_4
X_19691_ _23662_/Q VGND VGND VPWR VPWR _19691_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ _18642_/A _18636_/X _18639_/X _18641_/X VGND VGND VPWR VPWR _18642_/X sky130_fd_sc_hd__or4_4
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13407__A _13186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15854_ _15668_/B _15854_/B VGND VGND VPWR VPWR _15854_/X sky130_fd_sc_hd__or2_4
XFILLER_76_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14805_ scl_oen_o_S5 _14804_/Y _23985_/Q VGND VGND VPWR VPWR _14816_/B sky130_fd_sc_hd__and3_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18573_ _18479_/D _18573_/B VGND VGND VPWR VPWR _18573_/X sky130_fd_sc_hd__or2_4
X_15785_ _15561_/Y _15655_/X _15782_/X _21025_/B _15784_/X VGND VGND VPWR VPWR _15785_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12997_ _12323_/Y _12312_/X _12997_/C _12997_/D VGND VGND VPWR VPWR _12998_/C sky130_fd_sc_hd__or4_4
XFILLER_92_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19375__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17524_ _17517_/X _17524_/B _17521_/X _17524_/D VGND VGND VPWR VPWR _17524_/X sky130_fd_sc_hd__or4_4
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14736_ _22055_/A VGND VGND VPWR VPWR _14736_/Y sky130_fd_sc_hd__inv_2
X_11948_ _19632_/A VGND VGND VPWR VPWR _11948_/X sky130_fd_sc_hd__buf_2
XFILLER_60_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17455_ _13606_/X VGND VGND VPWR VPWR _17455_/X sky130_fd_sc_hd__buf_2
X_14667_ _14667_/A _13628_/X VGND VGND VPWR VPWR _14798_/A sky130_fd_sc_hd__or2_4
X_11879_ _11879_/A VGND VGND VPWR VPWR _17711_/A sky130_fd_sc_hd__inv_2
XANTENNA__24489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19127__B1 _19012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _16405_/Y _16403_/X _16315_/X _16403_/X VGND VGND VPWR VPWR _24608_/D sky130_fd_sc_hd__a2bb2o_4
X_13618_ _19346_/B _13617_/Y VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__and2_4
X_17386_ _17389_/A _17389_/B VGND VGND VPWR VPWR _17390_/B sky130_fd_sc_hd__or2_4
X_14598_ _25098_/Q _14578_/Y VGND VGND VPWR VPWR _14598_/X sky130_fd_sc_hd__or2_4
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19125_ _13272_/B VGND VGND VPWR VPWR _19125_/Y sky130_fd_sc_hd__inv_2
X_16337_ _16336_/Y _16333_/X _16238_/X _16333_/X VGND VGND VPWR VPWR _24632_/D sky130_fd_sc_hd__a2bb2o_4
X_13549_ _15701_/A _15920_/B VGND VGND VPWR VPWR _13601_/A sky130_fd_sc_hd__or2_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19056_ _19061_/A VGND VGND VPWR VPWR _19056_/X sky130_fd_sc_hd__buf_2
X_16268_ _16268_/A VGND VGND VPWR VPWR _16268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18007_ _18090_/A _19034_/A VGND VGND VPWR VPWR _18010_/B sky130_fd_sc_hd__or2_4
XANTENNA__21237__A1 _21046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15219_ _15243_/A _15053_/X _15218_/X VGND VGND VPWR VPWR _15219_/X sky130_fd_sc_hd__or3_4
XANTENNA__22434__B1 _22431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _23309_/A VGND VGND VPWR VPWR _16199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14911__B2 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22902__B _15681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12922__B1 _12875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23286__A _23263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19958_ _19958_/A VGND VGND VPWR VPWR _19958_/X sky130_fd_sc_hd__buf_2
XFILLER_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_108_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18909_ _18904_/Y _18907_/X _18908_/X _18907_/X VGND VGND VPWR VPWR _23934_/D sky130_fd_sc_hd__a2bb2o_4
X_19889_ _22026_/B _19883_/X _19632_/X _19888_/X VGND VGND VPWR VPWR _23594_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21920_ _21916_/X _21919_/X _22214_/A VGND VGND VPWR VPWR _21920_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21851_ _21848_/X _21851_/B _21850_/X VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__and3_4
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20802_ _13145_/B _13144_/X _20801_/Y VGND VGND VPWR VPWR _20802_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19004__A _19020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21782_ _22388_/A _21782_/B VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__or2_4
X_24570_ _24537_/CLK _24570_/D HRESETn VGND VGND VPWR VPWR _24570_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _25491_/CLK _20089_/X VGND VGND VPWR VPWR _13321_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_212_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20733_ _15625_/Y _20716_/X _20724_/X _20732_/Y VGND VGND VPWR VPWR _20734_/A sky130_fd_sc_hd__o22a_4
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24841__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _17405_/A _20661_/A VGND VGND VPWR VPWR _20664_/Y sky130_fd_sc_hd__nand2_4
X_23452_ _24684_/CLK _20280_/X VGND VGND VPWR VPWR _20276_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_46_0_HCLK clkbuf_8_46_0_HCLK/A VGND VGND VPWR VPWR _23690_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15942__A3 _15562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22403_ _23692_/Q _20344_/X VGND VGND VPWR VPWR _22403_/X sky130_fd_sc_hd__or2_4
XANTENNA__20180__A2_N _20177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23383_ _21026_/X VGND VGND VPWR VPWR IRQ[27] sky130_fd_sc_hd__buf_2
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17459__A _17459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20595_ _20594_/X VGND VGND VPWR VPWR _23958_/D sky130_fd_sc_hd__inv_2
XFILLER_164_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25122_ _25125_/CLK _14495_/X HRESETn VGND VGND VPWR VPWR _14494_/A sky130_fd_sc_hd__dfrtp_4
X_22334_ _15470_/Y _22334_/B VGND VGND VPWR VPWR _22334_/Y sky130_fd_sc_hd__nor2_4
XFILLER_192_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22265_ _22265_/A _22265_/B _22265_/C VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__and3_4
X_25053_ _24340_/CLK _14863_/X HRESETn VGND VGND VPWR VPWR _14824_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21216_ _20360_/A _21380_/A VGND VGND VPWR VPWR _21216_/X sky130_fd_sc_hd__or2_4
X_24004_ _24003_/CLK _24004_/D HRESETn VGND VGND VPWR VPWR _24004_/Q sky130_fd_sc_hd__dfrtp_4
X_22196_ _22190_/X _22192_/Y _22194_/Y _22195_/X _21565_/Y VGND VGND VPWR VPWR _22196_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_132_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21147_ _25308_/Q _12102_/X _13474_/Y _12102_/X VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21078_ _25525_/Q _21067_/X _21068_/X _21077_/X VGND VGND VPWR VPWR _21078_/X sky130_fd_sc_hd__a211o_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12920_ _12920_/A VGND VGND VPWR VPWR _25393_/D sky130_fd_sc_hd__inv_2
X_20029_ _20016_/Y VGND VGND VPWR VPWR _20029_/X sky130_fd_sc_hd__buf_2
X_24906_ _24493_/CLK _15627_/X HRESETn VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12851_ _12851_/A _12952_/C _12828_/A _12770_/Y VGND VGND VPWR VPWR _12856_/C sky130_fd_sc_hd__or4_4
X_24837_ _24883_/CLK _15832_/X HRESETn VGND VGND VPWR VPWR _24837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11802_/A VGND VGND VPWR VPWR _11802_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15589_/A VGND VGND VPWR VPWR _15626_/A sky130_fd_sc_hd__buf_2
XPHY_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _25397_/Q _24814_/Q _12780_/Y _12781_/Y VGND VGND VPWR VPWR _12786_/C sky130_fd_sc_hd__o22a_4
X_24768_ _24765_/CLK _24768_/D HRESETn VGND VGND VPWR VPWR _22758_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14510_/B VGND VGND VPWR VPWR _14521_/Y sky130_fd_sc_hd__inv_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _12077_/A _11733_/B VGND VGND VPWR VPWR _11734_/B sky130_fd_sc_hd__or2_4
X_23719_ _23678_/CLK _23719_/D VGND VGND VPWR VPWR _23719_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15918__B1 _24790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24699_ _24689_/CLK _16144_/X HRESETn VGND VGND VPWR VPWR _22673_/A sky130_fd_sc_hd__dfrtp_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24582__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17240_/A _17240_/B VGND VGND VPWR VPWR _17240_/X sky130_fd_sc_hd__or2_4
XFILLER_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14450_/Y _14446_/X _14427_/X _14451_/X VGND VGND VPWR VPWR _25140_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A VGND VGND VPWR VPWR _11710_/B sky130_fd_sc_hd__inv_2
XFILLER_187_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13371_/A _13403_/B VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__or2_4
XFILLER_186_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _17002_/A _17170_/Y VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__or2_4
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _14382_/Y VGND VGND VPWR VPWR _20463_/A sky130_fd_sc_hd__buf_2
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _22994_/A VGND VGND VPWR VPWR _16122_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13369_/A _19750_/A VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__or2_4
XFILLER_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16053_ _16053_/A VGND VGND VPWR VPWR _16053_/Y sky130_fd_sc_hd__inv_2
X_13265_ _13187_/X _13253_/X _13264_/X VGND VGND VPWR VPWR _13265_/X sky130_fd_sc_hd__and3_4
X_15004_ _15182_/B _24479_/Q _15003_/A _24479_/Q VGND VGND VPWR VPWR _15004_/X sky130_fd_sc_hd__a2bb2o_4
X_12216_ _24777_/Q VGND VGND VPWR VPWR _12216_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ _13199_/A _18958_/A VGND VGND VPWR VPWR _13197_/C sky130_fd_sc_hd__or2_4
XANTENNA__15817__A1_N _12377_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19812_ _19812_/A VGND VGND VPWR VPWR _21247_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _24115_/Q _12135_/B _12146_/Y VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__o21a_4
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19743_ _19742_/Y VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12078_ _13798_/B _21031_/A VGND VGND VPWR VPWR _21580_/A sky130_fd_sc_hd__or2_4
X_16955_ _16169_/Y _24266_/Q _21444_/A _16936_/X VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15906_ _12764_/Y _15904_/X _15905_/X _15904_/X VGND VGND VPWR VPWR _24800_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17832__A _17832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16886_ _16884_/Y _16877_/X _16885_/X _16877_/X VGND VGND VPWR VPWR _24414_/D sky130_fd_sc_hd__a2bb2o_4
X_19674_ _18334_/X _19075_/B _18938_/C VGND VGND VPWR VPWR _19675_/A sky130_fd_sc_hd__or3_4
XFILLER_225_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15837_ _12340_/Y _15835_/X _15765_/X _15835_/X VGND VGND VPWR VPWR _15837_/X sky130_fd_sc_hd__a2bb2o_4
X_18625_ _24538_/Q _24149_/Q _16586_/Y _18765_/A VGND VGND VPWR VPWR _18632_/A sky130_fd_sc_hd__o22a_4
XANTENNA__14458__A1_N _14178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16448__A _24588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15768_ _15772_/A VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__buf_2
X_18556_ _18493_/A VGND VGND VPWR VPWR _18556_/X sky130_fd_sc_hd__buf_2
XANTENNA__17270__C _17270_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14719_ _25068_/Q VGND VGND VPWR VPWR _14719_/Y sky130_fd_sc_hd__inv_2
X_17507_ _17507_/A _17503_/X _17507_/C _17506_/X VGND VGND VPWR VPWR _17507_/X sky130_fd_sc_hd__or4_4
X_18487_ _18487_/A _18486_/X VGND VGND VPWR VPWR _18487_/X sky130_fd_sc_hd__or2_4
XANTENNA__15909__B1 _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15699_ _15696_/B _15696_/C VGND VGND VPWR VPWR _15699_/X sky130_fd_sc_hd__or2_4
XFILLER_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17438_ _24334_/Q VGND VGND VPWR VPWR _21733_/A sky130_fd_sc_hd__inv_2
XFILLER_178_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16582__B1 _16412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_5_0_HCLK clkbuf_7_2_0_HCLK/X VGND VGND VPWR VPWR _23717_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_221_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17369_ _24355_/Q _17369_/B VGND VGND VPWR VPWR _17371_/B sky130_fd_sc_hd__or2_4
XANTENNA__22655__B1 _21844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19108_ _21906_/B _19105_/X _16885_/X _19105_/X VGND VGND VPWR VPWR _23865_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20380_ _21480_/B _20377_/X _19646_/A _20377_/X VGND VGND VPWR VPWR _23413_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22670__A3 _21550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14415__B _14388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19039_ _18090_/B VGND VGND VPWR VPWR _19039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22050_ _21499_/X _22049_/X _17738_/A VGND VGND VPWR VPWR _22050_/Y sky130_fd_sc_hd__a21oi_4
X_21001_ sda_oen_o_S4 _25104_/Q _20996_/A _14047_/A _21000_/Y VGND VGND VPWR VPWR
+ _23941_/D sky130_fd_sc_hd__a32o_4
XFILLER_217_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22952_ _22923_/X _22930_/X _22936_/Y _22951_/X VGND VGND VPWR VPWR HRDATA[19] sky130_fd_sc_hd__a211o_4
XFILLER_83_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21903_ _21412_/A VGND VGND VPWR VPWR _22380_/A sky130_fd_sc_hd__buf_2
XANTENNA__21264__A _21267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22883_ _22883_/A _22882_/X VGND VGND VPWR VPWR _22883_/X sky130_fd_sc_hd__or2_4
XANTENNA__12886__A _12638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19339__B1 _19226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16358__A _24623_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11790__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24622_ _24625_/CLK _16362_/X HRESETn VGND VGND VPWR VPWR _24622_/Q sky130_fd_sc_hd__dfrtp_4
X_21834_ _21834_/A _21660_/X VGND VGND VPWR VPWR _21839_/B sky130_fd_sc_hd__or2_4
XFILLER_243_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24553_ _24556_/CLK _24553_/D HRESETn VGND VGND VPWR VPWR _24553_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21765_ _21611_/X _21763_/X _21764_/X VGND VGND VPWR VPWR _21765_/X sky130_fd_sc_hd__and3_4
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23504_ _23488_/CLK _23504_/D VGND VGND VPWR VPWR _23504_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20716_ _20716_/A VGND VGND VPWR VPWR _20716_/X sky130_fd_sc_hd__buf_2
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24484_ _24485_/CLK _24484_/D HRESETn VGND VGND VPWR VPWR _24484_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16573__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21696_ _21815_/A _21694_/X _21696_/C VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__and3_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15915__A3 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _23555_/CLK _23435_/D VGND VGND VPWR VPWR _23435_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20647_ _17401_/A _17400_/X VGND VGND VPWR VPWR _20648_/B sky130_fd_sc_hd__nand2_4
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22110__A2 _22299_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20578_ _20578_/A VGND VGND VPWR VPWR _23954_/D sky130_fd_sc_hd__inv_2
X_23366_ VGND VGND VPWR VPWR _23366_/HI IRQ[30] sky130_fd_sc_hd__conb_1
XANTENNA__22823__A _22944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25105_ _25105_/CLK _14558_/X HRESETn VGND VGND VPWR VPWR sda_oen_o_S4 sky130_fd_sc_hd__dfstp_4
XANTENNA__23975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22317_ _24458_/Q _21312_/B _21335_/X VGND VGND VPWR VPWR _22317_/X sky130_fd_sc_hd__o21a_4
X_23297_ _22563_/X _23296_/X _22145_/C _11754_/A _23129_/X VGND VGND VPWR VPWR _23297_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13050_ _13049_/X VGND VGND VPWR VPWR _25362_/D sky130_fd_sc_hd__inv_2
X_25036_ _25043_/CLK _25036_/D HRESETn VGND VGND VPWR VPWR _14964_/A sky130_fd_sc_hd__dfrtp_4
X_22248_ _18314_/X VGND VGND VPWR VPWR _22264_/A sky130_fd_sc_hd__buf_2
XANTENNA__25128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12001_ _24105_/Q _12000_/X VGND VGND VPWR VPWR _12001_/X sky130_fd_sc_hd__and2_4
XFILLER_79_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12362__B2 _24838_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22179_ _22179_/A VGND VGND VPWR VPWR _22179_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16740_ _16736_/Y _16739_/X _16385_/X _16739_/X VGND VGND VPWR VPWR _16740_/X sky130_fd_sc_hd__a2bb2o_4
X_13952_ _13944_/A _13950_/Y _13952_/C _13952_/D VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__or4_4
XFILLER_247_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12903_ _12902_/X VGND VGND VPWR VPWR _12903_/Y sky130_fd_sc_hd__inv_2
X_16671_ _16671_/A VGND VGND VPWR VPWR _16671_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18250__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13883_ _21847_/A _13870_/X _25252_/Q _13872_/X VGND VGND VPWR VPWR _13883_/X sky130_fd_sc_hd__o22a_4
XFILLER_207_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12796__A _25375_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24763__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15622_ _22577_/A _15621_/X _11831_/X _15621_/X VGND VGND VPWR VPWR _24908_/D sky130_fd_sc_hd__a2bb2o_4
X_18410_ _16278_/Y _24163_/Q _16278_/Y _24163_/Q VGND VGND VPWR VPWR _18411_/D sky130_fd_sc_hd__a2bb2o_4
X_12834_ _25393_/Q VGND VGND VPWR VPWR _12834_/Y sky130_fd_sc_hd__inv_2
X_19390_ _19143_/A _19143_/B _19054_/C _19054_/D VGND VGND VPWR VPWR _19391_/A sky130_fd_sc_hd__and4_4
XANTENNA__16800__B2 _16738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18341_ _17477_/B _17459_/A VGND VGND VPWR VPWR _18342_/A sky130_fd_sc_hd__or2_4
X_15553_ _22575_/A VGND VGND VPWR VPWR _15553_/X sky130_fd_sc_hd__buf_2
X_12765_ _25399_/Q VGND VGND VPWR VPWR _12765_/Y sky130_fd_sc_hd__inv_2
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _20613_/A VGND VGND VPWR VPWR _14504_/X sky130_fd_sc_hd__buf_2
XANTENNA__22717__B _21855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _14684_/A VGND VGND VPWR VPWR _11718_/A sky130_fd_sc_hd__inv_2
X_18272_ _13804_/D _18262_/X _15993_/X _24229_/Q _18269_/X VGND VGND VPWR VPWR _18272_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_159_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15482_/Y _15477_/X _15483_/X _15477_/X VGND VGND VPWR VPWR _15484_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12683_/X VGND VGND VPWR VPWR _12697_/B sky130_fd_sc_hd__inv_2
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17223_ _16329_/Y _17212_/A _24638_/Q _17322_/A VGND VGND VPWR VPWR _17223_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _14428_/A VGND VGND VPWR VPWR _14435_/X sky130_fd_sc_hd__buf_2
XANTENNA__17099__A _17064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13420__A _13420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _17127_/X _17142_/B _17153_/Y VGND VGND VPWR VPWR _17154_/X sky130_fd_sc_hd__and3_4
XFILLER_168_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14366_ MSO_S3 _14365_/X _25165_/Q _14360_/X VGND VGND VPWR VPWR _14366_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__16316__B1 _16315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_92_0_HCLK clkbuf_7_46_0_HCLK/X VGND VGND VPWR VPWR _24878_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_183_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16105_ _16102_/Y _16098_/X _15948_/X _16104_/X VGND VGND VPWR VPWR _24715_/D sky130_fd_sc_hd__a2bb2o_4
X_13317_ _13317_/A _23913_/Q VGND VGND VPWR VPWR _13318_/C sky130_fd_sc_hd__or2_4
X_17085_ _17084_/X VGND VGND VPWR VPWR _17085_/Y sky130_fd_sc_hd__inv_2
X_14297_ _14309_/A VGND VGND VPWR VPWR _14305_/A sky130_fd_sc_hd__inv_2
XFILLER_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25551__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16731__A _16379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16036_ _16019_/A VGND VGND VPWR VPWR _16036_/X sky130_fd_sc_hd__buf_2
XFILLER_182_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13248_ _13155_/X VGND VGND VPWR VPWR _13249_/A sky130_fd_sc_hd__buf_2
XANTENNA__11875__A _13818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _13198_/A _13179_/B VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__or2_4
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13793__C _13804_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17987_ _17987_/A _17987_/B VGND VGND VPWR VPWR _17988_/C sky130_fd_sc_hd__or2_4
XANTENNA__19569__B1 _19454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19726_ _19724_/Y _19720_/X _19659_/X _19725_/X VGND VGND VPWR VPWR _19726_/X sky130_fd_sc_hd__a2bb2o_4
X_16938_ _21444_/A _16936_/X _22162_/A _16937_/Y VGND VGND VPWR VPWR _16941_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19657_ _19655_/Y _19653_/X _19656_/X _19653_/X VGND VGND VPWR VPWR _19657_/X sky130_fd_sc_hd__a2bb2o_4
X_16869_ _16867_/Y _16868_/X RsRx_S0 _16868_/X VGND VGND VPWR VPWR _16869_/X sky130_fd_sc_hd__a2bb2o_4
X_18608_ _24137_/Q VGND VGND VPWR VPWR _18691_/B sky130_fd_sc_hd__inv_2
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19588_ _21694_/B _19587_/X _11961_/X _19587_/X VGND VGND VPWR VPWR _19588_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18539_ _18539_/A _18539_/B VGND VGND VPWR VPWR _18543_/B sky130_fd_sc_hd__or2_4
XFILLER_240_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21550_ _21314_/A VGND VGND VPWR VPWR _21550_/X sky130_fd_sc_hd__buf_2
XFILLER_221_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21531__B _23016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16555__B1 _16385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20501_ _20537_/A _20501_/B VGND VGND VPWR VPWR _24091_/D sky130_fd_sc_hd__or2_4
X_21481_ _21676_/A _20031_/Y VGND VGND VPWR VPWR _21481_/X sky130_fd_sc_hd__or2_4
XFILLER_166_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14426__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20432_ _13353_/B VGND VGND VPWR VPWR _20432_/Y sky130_fd_sc_hd__inv_2
X_23220_ _16564_/A _22485_/X _22852_/X _23219_/X VGND VGND VPWR VPWR _23221_/C sky130_fd_sc_hd__a211o_4
XFILLER_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16307__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20363_ _19965_/A _19480_/X _19481_/X VGND VGND VPWR VPWR _20364_/A sky130_fd_sc_hd__or3_4
X_23151_ _23013_/A _23147_/X _23151_/C VGND VGND VPWR VPWR _23151_/X sky130_fd_sc_hd__and3_4
XANTENNA__25292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_0_0_HCLK clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_173_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22102_ _15135_/A _23274_/B VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__or2_4
X_23082_ _16822_/A _22947_/X _23015_/X _23081_/X VGND VGND VPWR VPWR _23082_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14333__A2 _25175_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20294_ _21414_/B _20291_/X _19810_/A _20291_/X VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22033_ _22029_/A _22033_/B _22032_/X VGND VGND VPWR VPWR _22033_/X sky130_fd_sc_hd__and3_4
XANTENNA__21603__A1 _21606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23193__B _23189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23984_ _24003_/CLK _23984_/D HRESETn VGND VGND VPWR VPWR _23984_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22935_ _22801_/X _22932_/X _22804_/X _22934_/X VGND VGND VPWR VPWR _22936_/B sky130_fd_sc_hd__o22a_4
XFILLER_217_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19980__B1 _19643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22866_ _22771_/X _22863_/X _22446_/A _22865_/X VGND VGND VPWR VPWR _22866_/X sky130_fd_sc_hd__o22a_4
XFILLER_204_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24605_ _24602_/CLK _24605_/D HRESETn VGND VGND VPWR VPWR _24605_/Q sky130_fd_sc_hd__dfrtp_4
X_21817_ _21679_/A _21809_/X _21817_/C VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__or3_4
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22797_ _12197_/X _22507_/X _17767_/A _21079_/A VGND VGND VPWR VPWR _22799_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16816__A _16810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ _12550_/A VGND VGND VPWR VPWR _12550_/Y sky130_fd_sc_hd__inv_2
X_24536_ _24601_/CLK _24536_/D HRESETn VGND VGND VPWR VPWR _24536_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21748_ _22941_/A VGND VGND VPWR VPWR _22542_/A sky130_fd_sc_hd__buf_2
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13544__A1_N SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22619__B1 _21844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12229_/X _12212_/X _12288_/Y _12480_/X VGND VGND VPWR VPWR _12481_/X sky130_fd_sc_hd__or4_4
X_24467_ _24430_/CLK _24467_/D HRESETn VGND VGND VPWR VPWR _15012_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21679_ _21679_/A _21671_/X _21678_/X VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__or3_4
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _14218_/Y _14219_/X _13812_/X _14210_/X VGND VGND VPWR VPWR _14220_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23418_ _23563_/CLK _20368_/X VGND VGND VPWR VPWR _23418_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _24240_/CLK _17108_/Y HRESETn VGND VGND VPWR VPWR _24398_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_79_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14151_ _14111_/A _14111_/B _14111_/A _14111_/B VGND VGND VPWR VPWR _14151_/X sky130_fd_sc_hd__a2bb2o_4
X_23349_ _22813_/A _23340_/Y _23349_/C _23348_/X VGND VGND VPWR VPWR _23349_/X sky130_fd_sc_hd__or4_4
XANTENNA__16551__A _15718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _13104_/A _13102_/B _13102_/C VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__and3_4
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14082_ _14082_/A _14082_/B VGND VGND VPWR VPWR _14082_/X sky130_fd_sc_hd__and2_4
XANTENNA__12185__A1_N _14338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23044__B1 _11782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23087__C _22954_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13033_ _13044_/A _13031_/X _13032_/X VGND VGND VPWR VPWR _25367_/D sky130_fd_sc_hd__and3_4
X_17910_ _17900_/Y _17910_/B VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__and2_4
X_25019_ _25018_/CLK _25019_/D HRESETn VGND VGND VPWR VPWR _25019_/Q sky130_fd_sc_hd__dfrtp_4
X_18890_ _18890_/A VGND VGND VPWR VPWR _18890_/X sky130_fd_sc_hd__buf_2
XFILLER_154_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17841_ _17843_/B VGND VGND VPWR VPWR _17842_/B sky130_fd_sc_hd__inv_2
XFILLER_79_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14984_ _14984_/A VGND VGND VPWR VPWR _14990_/A sky130_fd_sc_hd__inv_2
X_17772_ _17750_/Y _17771_/X VGND VGND VPWR VPWR _17793_/B sky130_fd_sc_hd__or2_4
XFILLER_207_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19511_ _22267_/B _19508_/X _11943_/X _19508_/X VGND VGND VPWR VPWR _23723_/D sky130_fd_sc_hd__a2bb2o_4
X_13935_ _24979_/Q _13933_/X _13942_/A _13934_/X VGND VGND VPWR VPWR _13935_/X sky130_fd_sc_hd__or4_4
X_16723_ _16723_/A VGND VGND VPWR VPWR _16723_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16654_ _16709_/A VGND VGND VPWR VPWR _16654_/X sky130_fd_sc_hd__buf_2
X_19442_ _19441_/Y _19438_/X _19418_/X _19438_/X VGND VGND VPWR VPWR _23747_/D sky130_fd_sc_hd__a2bb2o_4
X_13866_ _13864_/X _13876_/A _13871_/A VGND VGND VPWR VPWR _13866_/X sky130_fd_sc_hd__a21o_4
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22728__A _21714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15605_ _15604_/Y _15602_/X _11800_/X _15602_/X VGND VGND VPWR VPWR _24915_/D sky130_fd_sc_hd__a2bb2o_4
X_12817_ _12817_/A VGND VGND VPWR VPWR _12817_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21632__A _14709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16585_ _16583_/Y _16579_/X _16414_/X _16584_/X VGND VGND VPWR VPWR _16585_/X sky130_fd_sc_hd__a2bb2o_4
X_19373_ _23770_/Q VGND VGND VPWR VPWR _19373_/Y sky130_fd_sc_hd__inv_2
X_13797_ _11733_/B VGND VGND VPWR VPWR _17448_/B sky130_fd_sc_hd__buf_2
XANTENNA__16726__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15050__A1_N _25019_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15536_ _15653_/A _15533_/X HADDR[8] _15533_/X VGND VGND VPWR VPWR _24938_/D sky130_fd_sc_hd__a2bb2o_4
X_18324_ _20015_/B _18323_/X _18286_/Y _18323_/X VGND VGND VPWR VPWR _18324_/X sky130_fd_sc_hd__a2bb2o_4
X_12748_ _12747_/X VGND VGND VPWR VPWR _12748_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21323__A2_N _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18255_ _18245_/X _18247_/X _16609_/X _22525_/A _18248_/X VGND VGND VPWR VPWR _18255_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15467_ _14289_/X _14260_/A _15440_/X _13927_/B _15461_/X VGND VGND VPWR VPWR _15467_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12679_ _12679_/A _12676_/X VGND VGND VPWR VPWR _12680_/C sky130_fd_sc_hd__or2_4
XANTENNA__16439__A1_N _15121_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _17205_/Y VGND VGND VPWR VPWR _17364_/A sky130_fd_sc_hd__buf_2
X_14418_ _14428_/A VGND VGND VPWR VPWR _14418_/X sky130_fd_sc_hd__buf_2
X_18186_ _17975_/X _18184_/X _18186_/C VGND VGND VPWR VPWR _18186_/X sky130_fd_sc_hd__and3_4
XFILLER_128_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15398_ _15153_/Y _15397_/X VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__or2_4
XFILLER_156_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17137_ _17048_/Y _17137_/B _17053_/C _17136_/X VGND VGND VPWR VPWR _17138_/B sky130_fd_sc_hd__or4_4
X_14349_ _14349_/A _14347_/Y _14349_/C _14349_/D VGND VGND VPWR VPWR _14350_/A sky130_fd_sc_hd__or4_4
XFILLER_144_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16461__A _22944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17068_ _17074_/A _17068_/B VGND VGND VPWR VPWR _17079_/A sky130_fd_sc_hd__or2_4
XANTENNA__21079__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16019_ _16019_/A VGND VGND VPWR VPWR _16019_/X sky130_fd_sc_hd__buf_2
XANTENNA__19772__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24685__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24614__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19709_ _19708_/Y _19704_/X _19612_/X _19704_/X VGND VGND VPWR VPWR _23656_/D sky130_fd_sc_hd__a2bb2o_4
X_20981_ _20981_/A _20982_/B VGND VGND VPWR VPWR _20981_/X sky130_fd_sc_hd__and2_4
XFILLER_226_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22720_ _24360_/Q _21868_/B VGND VGND VPWR VPWR _22723_/B sky130_fd_sc_hd__or2_4
XFILLER_92_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22651_ _22651_/A _22577_/B VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__and2_4
XFILLER_81_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22313__A2 _21450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21602_ _15643_/Y _21330_/A VGND VGND VPWR VPWR _21602_/X sky130_fd_sc_hd__and2_4
XANTENNA__19012__A _19151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15540__A _21135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25370_ _25365_/CLK _25370_/D HRESETn VGND VGND VPWR VPWR _25370_/Q sky130_fd_sc_hd__dfrtp_4
X_22582_ _22582_/A VGND VGND VPWR VPWR _22582_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16528__B1 _16157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24321_ _23534_/CLK _24321_/D HRESETn VGND VGND VPWR VPWR _17572_/A sky130_fd_sc_hd__dfrtp_4
X_21533_ _21530_/X _21531_/X _21532_/X _25527_/Q _22530_/B VGND VGND VPWR VPWR _21533_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24252_ _24252_/CLK _18071_/X HRESETn VGND VGND VPWR VPWR _24252_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21464_ _17716_/A VGND VGND VPWR VPWR _21815_/A sky130_fd_sc_hd__buf_2
XFILLER_147_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22373__A _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23203_ _23124_/X _23202_/X _23058_/X _24748_/Q _22990_/X VGND VGND VPWR VPWR _23203_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_181_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20415_ _20408_/X _20404_/X _15993_/X _23399_/Q _20406_/X VGND VGND VPWR VPWR _23399_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_146_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21395_ _21246_/A _21393_/X _21394_/X VGND VGND VPWR VPWR _21395_/X sky130_fd_sc_hd__and3_4
X_24183_ _24189_/CLK _24183_/D HRESETn VGND VGND VPWR VPWR _24183_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23134_ _17305_/A _22926_/X _12899_/A _22927_/X VGND VGND VPWR VPWR _23134_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20346_ _20345_/X VGND VGND VPWR VPWR _20346_/X sky130_fd_sc_hd__buf_2
XANTENNA__16700__B1 _15759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19682__A _19675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20277_ _19859_/X _20149_/B _19278_/X VGND VGND VPWR VPWR _20278_/A sky130_fd_sc_hd__or3_4
X_23065_ _23208_/A _23065_/B _23065_/C _23064_/X VGND VGND VPWR VPWR _23065_/X sky130_fd_sc_hd__or4_4
XFILLER_68_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22820__B _15681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22016_ _20410_/Y _22013_/Y _22014_/X _22015_/Y VGND VGND VPWR VPWR _22017_/A sky130_fd_sc_hd__a211o_4
XANTENNA__23329__A1 _22563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23329__B2 _22565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15715__A _21172_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22537__C1 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11828__B1 _11827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11981_ _11970_/C _11712_/A VGND VGND VPWR VPWR _11981_/X sky130_fd_sc_hd__or2_4
X_23967_ _24095_/CLK _23967_/D HRESETn VGND VGND VPWR VPWR _14543_/A sky130_fd_sc_hd__dfstp_4
XFILLER_17_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13720_ _13700_/B _13716_/X _13719_/Y _13712_/X _11688_/A VGND VGND VPWR VPWR _25296_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13235__A _13356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22918_ _22788_/X _22917_/X _22497_/X _24740_/Q _22498_/X VGND VGND VPWR VPWR _22919_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23898_ _23880_/CLK _23898_/D VGND VGND VPWR VPWR _23898_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22548__A _22592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21452__A _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13651_ _13649_/X _13650_/X VGND VGND VPWR VPWR _25306_/D sky130_fd_sc_hd__or2_4
XFILLER_204_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22849_ _22738_/A VGND VGND VPWR VPWR _22849_/X sky130_fd_sc_hd__buf_2
XFILLER_140_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12602_ _12601_/Y _24890_/Q _12601_/Y _24890_/Q VGND VGND VPWR VPWR _12602_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ _24619_/Q VGND VGND VPWR VPWR _16370_/Y sky130_fd_sc_hd__inv_2
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582_ _13582_/A VGND VGND VPWR VPWR _13582_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14793__A2 _14791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21512__B1 _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A _15321_/B VGND VGND VPWR VPWR _15323_/B sky130_fd_sc_hd__or2_4
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12533_ _25432_/Q VGND VGND VPWR VPWR _12630_/A sky130_fd_sc_hd__inv_2
X_24519_ _24684_/CLK _24519_/D HRESETn VGND VGND VPWR VPWR _13749_/A sky130_fd_sc_hd__dfrtp_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25499_ _24201_/CLK _25499_/D HRESETn VGND VGND VPWR VPWR _25499_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18040_ _17987_/A _23466_/Q VGND VGND VPWR VPWR _18040_/X sky130_fd_sc_hd__or2_4
XFILLER_173_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15252_ _15252_/A _15252_/B _15252_/C VGND VGND VPWR VPWR _15252_/X sky130_fd_sc_hd__and3_4
XFILLER_184_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12464_ _12464_/A _12464_/B VGND VGND VPWR VPWR _12465_/C sky130_fd_sc_hd__or2_4
XANTENNA__23379__A _21022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22283__A _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14203_ _14202_/X VGND VGND VPWR VPWR _14203_/X sky130_fd_sc_hd__buf_2
XFILLER_126_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12556__B2 _12555_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15183_ _14996_/A VGND VGND VPWR VPWR _15183_/X sky130_fd_sc_hd__buf_2
X_12395_ _12395_/A VGND VGND VPWR VPWR _12395_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_11_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14134_ _14153_/A VGND VGND VPWR VPWR _14134_/X sky130_fd_sc_hd__buf_2
XFILLER_125_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23017__B1 _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19991_ _22366_/B _19989_/X _19990_/X _19989_/X VGND VGND VPWR VPWR _23556_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_103_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24915_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_153_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14065_ _14064_/X VGND VGND VPWR VPWR _14066_/A sky130_fd_sc_hd__buf_2
X_18942_ _18942_/A VGND VGND VPWR VPWR _18942_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17722__A1_N _21485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_166_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23459_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12314__A _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_9_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13016_ _13049_/A VGND VGND VPWR VPWR _13019_/A sky130_fd_sc_hd__buf_2
X_18873_ _18830_/Y _18729_/X _18851_/X _18872_/X VGND VGND VPWR VPWR _18873_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17824_ _17824_/A _17824_/B VGND VGND VPWR VPWR _17825_/C sky130_fd_sc_hd__or2_4
XFILLER_239_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11819__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ _25030_/Q VGND VGND VPWR VPWR _15232_/A sky130_fd_sc_hd__inv_2
X_17755_ _24267_/Q VGND VGND VPWR VPWR _17757_/C sky130_fd_sc_hd__inv_2
XFILLER_82_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16706_ _16706_/A VGND VGND VPWR VPWR _16706_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17840__A _17766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13918_ _13908_/A _13910_/A _13915_/A _13955_/B VGND VGND VPWR VPWR _13937_/B sky130_fd_sc_hd__or4_4
X_14898_ _15178_/A _16803_/A _15178_/A _16803_/A VGND VGND VPWR VPWR _14898_/X sky130_fd_sc_hd__a2bb2o_4
X_17686_ _17518_/Y _17676_/X VGND VGND VPWR VPWR _17687_/C sky130_fd_sc_hd__nand2_4
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19425_ _19424_/Y _19422_/X _19377_/X _19422_/X VGND VGND VPWR VPWR _19425_/X sky130_fd_sc_hd__a2bb2o_4
X_13849_ _11851_/A VGND VGND VPWR VPWR _13849_/X sky130_fd_sc_hd__buf_2
X_16637_ _14779_/A _14776_/C _16633_/X _13749_/A _16636_/X VGND VGND VPWR VPWR _24519_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15360__A _15388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19356_ _19355_/Y _19353_/X _19220_/X _19353_/X VGND VGND VPWR VPWR _19356_/X sky130_fd_sc_hd__a2bb2o_4
X_16568_ _16566_/Y _16567_/X _16306_/X _16567_/X VGND VGND VPWR VPWR _24546_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12795__A1 _12793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18307_ _18297_/X VGND VGND VPWR VPWR _18310_/B sky130_fd_sc_hd__inv_2
XFILLER_148_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15519_ _24944_/Q VGND VGND VPWR VPWR _15519_/Y sky130_fd_sc_hd__inv_2
X_16499_ _24571_/Q VGND VGND VPWR VPWR _16499_/Y sky130_fd_sc_hd__inv_2
X_19287_ _22077_/B _19281_/X _16881_/X _19286_/X VGND VGND VPWR VPWR _19287_/X sky130_fd_sc_hd__a2bb2o_4
X_18238_ _13824_/X VGND VGND VPWR VPWR _21974_/A sky130_fd_sc_hd__buf_2
XANTENNA__15733__A1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23256__B1 _22815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18169_ _18169_/A _18169_/B _18168_/X VGND VGND VPWR VPWR _18170_/C sky130_fd_sc_hd__and3_4
XANTENNA__16191__A _16190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20200_ _23481_/Q VGND VGND VPWR VPWR _20200_/Y sky130_fd_sc_hd__inv_2
X_21180_ _22527_/A VGND VGND VPWR VPWR _21180_/X sky130_fd_sc_hd__buf_2
XANTENNA__24866__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20131_ _20131_/A VGND VGND VPWR VPWR _20131_/Y sky130_fd_sc_hd__inv_2
X_20062_ _23531_/Q VGND VGND VPWR VPWR _20062_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21537__A _21537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24870_ _24867_/CLK _24870_/D HRESETn VGND VGND VPWR VPWR _24870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19007__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23821_ _23830_/CLK _23821_/D VGND VGND VPWR VPWR _19230_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17750__A _24289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23752_ _23754_/CLK _23752_/D VGND VGND VPWR VPWR _18117_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_226_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20964_ _20964_/A VGND VGND VPWR VPWR _20964_/Y sky130_fd_sc_hd__inv_2
XFILLER_242_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16749__B1 _15732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _12247_/X _22732_/A _17766_/B _22702_/X VGND VGND VPWR VPWR _22703_/X sky130_fd_sc_hd__o22a_4
XFILLER_226_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _23563_/CLK _23683_/D VGND VGND VPWR VPWR _23683_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _24061_/Q VGND VGND VPWR VPWR _20895_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14224__B2 _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25422_ _25425_/CLK _12695_/X HRESETn VGND VGND VPWR VPWR _25422_/Q sky130_fd_sc_hd__dfrtp_4
X_22634_ _17258_/Y _22677_/B _22633_/Y VGND VGND VPWR VPWR _22634_/X sky130_fd_sc_hd__o21a_4
XFILLER_179_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25353_ _25365_/CLK _13085_/X HRESETn VGND VGND VPWR VPWR _13083_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22565_ _11747_/A VGND VGND VPWR VPWR _22565_/X sky130_fd_sc_hd__buf_2
XFILLER_110_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24304_ _24302_/CLK _17687_/X HRESETn VGND VGND VPWR VPWR _24304_/Q sky130_fd_sc_hd__dfrtp_4
X_21516_ _21384_/B _21515_/X VGND VGND VPWR VPWR _21517_/C sky130_fd_sc_hd__or2_4
X_25284_ _23690_/CLK _25284_/D HRESETn VGND VGND VPWR VPWR _25284_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15724__A1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22496_ _24626_/Q _22789_/B VGND VGND VPWR VPWR _22496_/X sky130_fd_sc_hd__or2_4
XFILLER_155_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24235_ _24238_/CLK _24235_/D HRESETn VGND VGND VPWR VPWR _24235_/Q sky130_fd_sc_hd__dfrtp_4
X_21447_ _15565_/X _21444_/X _21445_/X _11869_/A _22530_/B VGND VGND VPWR VPWR _21447_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_154_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ _25471_/Q VGND VGND VPWR VPWR SSn_S3 sky130_fd_sc_hd__inv_2
X_24166_ _24192_/CLK _24166_/D HRESETn VGND VGND VPWR VPWR _24166_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22470__A1 _12113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21378_ _21565_/A _21378_/B VGND VGND VPWR VPWR _21378_/Y sky130_fd_sc_hd__nor2_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15488__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20481__B1 _14550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23117_ _23117_/A _23116_/X VGND VGND VPWR VPWR _23132_/B sky130_fd_sc_hd__and2_4
X_20329_ _20323_/Y VGND VGND VPWR VPWR _20329_/X sky130_fd_sc_hd__buf_2
XFILLER_123_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24097_ _25106_/CLK _20476_/X HRESETn VGND VGND VPWR VPWR _20444_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18452__A1_N _16271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17536__A2_N _17578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_239_0_HCLK clkbuf_8_238_0_HCLK/A VGND VGND VPWR VPWR _25246_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14160__B1 _25143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23048_ _23025_/X _23029_/X _23048_/C _23047_/X VGND VGND VPWR VPWR HRDATA[22] sky130_fd_sc_hd__or4_4
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15870_ _15710_/X _15870_/B VGND VGND VPWR VPWR _15896_/A sky130_fd_sc_hd__or2_4
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14821_ _14812_/C VGND VGND VPWR VPWR _14828_/A sky130_fd_sc_hd__inv_2
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24999_ _24981_/CLK _24999_/D HRESETn VGND VGND VPWR VPWR _24999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21355__A1_N _14186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14752_ _14751_/Y _14732_/Y _22056_/A _14731_/X VGND VGND VPWR VPWR _25070_/D sky130_fd_sc_hd__o22a_4
X_17540_ _11820_/Y _17581_/A _11820_/Y _17581_/A VGND VGND VPWR VPWR _17540_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11964_ _19646_/A VGND VGND VPWR VPWR _11964_/X sky130_fd_sc_hd__buf_2
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13703_ _13703_/A _13703_/B VGND VGND VPWR VPWR _13703_/X sky130_fd_sc_hd__or2_4
XFILLER_72_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17471_ _17471_/A _17470_/X VGND VGND VPWR VPWR _17484_/C sky130_fd_sc_hd__or2_4
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14683_ _14683_/A VGND VGND VPWR VPWR _14730_/C sky130_fd_sc_hd__inv_2
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11895_ _11894_/X VGND VGND VPWR VPWR _11895_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16276__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19210_ _19028_/B _19054_/C _19054_/D _19054_/A VGND VGND VPWR VPWR _19210_/X sky130_fd_sc_hd__and4_4
X_13634_ _14667_/A VGND VGND VPWR VPWR _13634_/X sky130_fd_sc_hd__buf_2
X_16422_ _16390_/A VGND VGND VPWR VPWR _16442_/A sky130_fd_sc_hd__buf_2
XANTENNA__25324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16353_ _16351_/Y _16346_/X _16153_/X _16352_/X VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__a2bb2o_4
X_19141_ _19141_/A VGND VGND VPWR VPWR _19141_/Y sky130_fd_sc_hd__inv_2
X_13565_ _13564_/Y _25103_/Q _13564_/Y _25103_/Q VGND VGND VPWR VPWR _13565_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16730__A2_N _16654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _25002_/Q VGND VGND VPWR VPWR _15365_/A sky130_fd_sc_hd__inv_2
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12516_ _13051_/A VGND VGND VPWR VPWR _13049_/A sky130_fd_sc_hd__inv_2
X_19072_ _19072_/A VGND VGND VPWR VPWR _19072_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16284_ _15681_/X VGND VGND VPWR VPWR _16284_/X sky130_fd_sc_hd__buf_2
XFILLER_9_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23238__B1 _25553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13496_ _13495_/Y _13491_/X _11862_/X _13491_/X VGND VGND VPWR VPWR _25325_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17819__B _17766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _15231_/X VGND VGND VPWR VPWR _15235_/Y sky130_fd_sc_hd__inv_2
X_18023_ _18023_/A _19193_/A VGND VGND VPWR VPWR _18023_/X sky130_fd_sc_hd__or2_4
XFILLER_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ _12269_/Y _12442_/B _12411_/X _12444_/B VGND VGND VPWR VPWR _12447_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_49_0_HCLK clkbuf_5_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _25009_/Q _15154_/Y _15153_/Y _16445_/A VGND VGND VPWR VPWR _15166_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22461__A1 _15017_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ _25360_/Q VGND VGND VPWR VPWR _13054_/A sky130_fd_sc_hd__inv_2
X_14117_ _14117_/A VGND VGND VPWR VPWR _14117_/X sky130_fd_sc_hd__buf_2
X_15097_ _24991_/Q _15095_/Y _15096_/Y _24611_/Q VGND VGND VPWR VPWR _15097_/X sky130_fd_sc_hd__a2bb2o_4
X_19974_ _23561_/Q VGND VGND VPWR VPWR _19974_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14048_ _13984_/A _14021_/B VGND VGND VPWR VPWR _14048_/Y sky130_fd_sc_hd__nand2_4
X_18925_ _21909_/B _18922_/X _16885_/X _18922_/X VGND VGND VPWR VPWR _18925_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23275__C _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18856_ _18852_/X _18856_/B _18854_/X _18855_/X VGND VGND VPWR VPWR _18856_/X sky130_fd_sc_hd__or4_4
XFILLER_227_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17807_ _17753_/A _17807_/B VGND VGND VPWR VPWR _17807_/X sky130_fd_sc_hd__or2_4
Xclkbuf_4_4_0_HCLK clkbuf_3_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18787_ _18749_/A VGND VGND VPWR VPWR _18806_/A sky130_fd_sc_hd__buf_2
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15999_ _15999_/A VGND VGND VPWR VPWR _15999_/Y sky130_fd_sc_hd__inv_2
X_17738_ _17738_/A VGND VGND VPWR VPWR _21509_/A sky130_fd_sc_hd__buf_2
XFILLER_236_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17669_ _17581_/Y _17664_/B _17666_/B _17600_/X VGND VGND VPWR VPWR _17670_/A sky130_fd_sc_hd__a211o_4
XFILLER_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19408_ _19407_/Y _19405_/X _19341_/X _19405_/X VGND VGND VPWR VPWR _23758_/D sky130_fd_sc_hd__a2bb2o_4
X_20680_ _20680_/A _20679_/X VGND VGND VPWR VPWR _20680_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19339_ _19337_/Y _19338_/X _19226_/X _19338_/X VGND VGND VPWR VPWR _23783_/D sky130_fd_sc_hd__a2bb2o_4
X_22350_ _21941_/A _20362_/Y VGND VGND VPWR VPWR _22350_/X sky130_fd_sc_hd__or2_4
XFILLER_176_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21301_ _21300_/Y VGND VGND VPWR VPWR _22202_/C sky130_fd_sc_hd__buf_2
X_22281_ _22281_/A VGND VGND VPWR VPWR _22281_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14434__A _25145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24020_ _24020_/CLK _20720_/Y HRESETn VGND VGND VPWR VPWR _13136_/A sky130_fd_sc_hd__dfrtp_4
X_21232_ _16728_/Y _21877_/B VGND VGND VPWR VPWR _21238_/B sky130_fd_sc_hd__or2_4
XANTENNA__18656__B1 _16578_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17745__A _17710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21163_ _14250_/Y _14229_/A _17445_/Y _21373_/A VGND VGND VPWR VPWR _21164_/D sky130_fd_sc_hd__o22a_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20114_ _23512_/Q VGND VGND VPWR VPWR _21791_/B sky130_fd_sc_hd__inv_2
XANTENNA__21267__A _21267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21094_ _21093_/X VGND VGND VPWR VPWR _21094_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11793__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20045_ _20043_/Y _20039_/X _19996_/X _20044_/X VGND VGND VPWR VPWR _20045_/X sky130_fd_sc_hd__a2bb2o_4
X_24922_ _24042_/CLK _15587_/X HRESETn VGND VGND VPWR VPWR _15586_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_69_0_HCLK clkbuf_7_34_0_HCLK/X VGND VGND VPWR VPWR _25380_/CLK sky130_fd_sc_hd__clkbuf_1
X_24853_ _24878_/CLK _15810_/X HRESETn VGND VGND VPWR VPWR _24853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15642__B1 _15483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23804_ _23475_/CLK _23804_/D VGND VGND VPWR VPWR _23804_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24784_ _24803_/CLK _24784_/D HRESETn VGND VGND VPWR VPWR _24784_/Q sky130_fd_sc_hd__dfrtp_4
X_21996_ _21996_/A _22275_/A _21996_/C _23424_/Q VGND VGND VPWR VPWR _21996_/X sky130_fd_sc_hd__or4_4
XPHY_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23735_/CLK _23735_/D VGND VGND VPWR VPWR _18152_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_226_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _24073_/Q VGND VGND VPWR VPWR _20947_/Y sky130_fd_sc_hd__inv_2
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _24242_/Q VGND VGND VPWR VPWR _22595_/A sky130_fd_sc_hd__inv_2
X_23666_ _23642_/CLK _23666_/D VGND VGND VPWR VPWR _19681_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_187_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20836_/A VGND VGND VPWR VPWR _20878_/X sky130_fd_sc_hd__buf_2
XFILLER_230_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22826__A _22944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25405_ _24824_/CLK _12750_/X HRESETn VGND VGND VPWR VPWR _21023_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22617_ _21123_/A _22615_/X _22121_/X _22616_/X VGND VGND VPWR VPWR _22618_/B sky130_fd_sc_hd__o22a_4
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23597_ _23597_/CLK _23597_/D VGND VGND VPWR VPWR _19878_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22140__B1 _12572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13350_ _13222_/X _13350_/B VGND VGND VPWR VPWR _13351_/C sky130_fd_sc_hd__or2_4
X_25336_ _25488_/CLK _25336_/D HRESETn VGND VGND VPWR VPWR _25336_/Q sky130_fd_sc_hd__dfrtp_4
X_22548_ _22592_/A _22548_/B _22547_/X VGND VGND VPWR VPWR _22548_/X sky130_fd_sc_hd__and3_4
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12301_ _12301_/A VGND VGND VPWR VPWR _13002_/C sky130_fd_sc_hd__inv_2
XANTENNA__24788__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13281_ _13356_/A _18944_/A VGND VGND VPWR VPWR _13283_/B sky130_fd_sc_hd__or2_4
X_25267_ _24230_/CLK _25267_/D HRESETn VGND VGND VPWR VPWR _13566_/A sky130_fd_sc_hd__dfrtp_4
X_22479_ _22479_/A _22479_/B VGND VGND VPWR VPWR _22480_/D sky130_fd_sc_hd__nor2_4
XFILLER_108_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15020_ _25015_/Q _15019_/A _15290_/A _15019_/Y VGND VGND VPWR VPWR _15021_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24717__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12232_ _25440_/Q VGND VGND VPWR VPWR _12232_/Y sky130_fd_sc_hd__inv_2
X_24218_ _24217_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _17714_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25198_ _24979_/CLK _14262_/X HRESETn VGND VGND VPWR VPWR sda_oen_o_S5 sky130_fd_sc_hd__dfstp_4
XANTENNA_clkbuf_5_3_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12163_ _24120_/Q _12162_/A _12161_/Y _12162_/Y VGND VGND VPWR VPWR _24120_/D sky130_fd_sc_hd__o22a_4
X_24149_ _24989_/CLK _24149_/D HRESETn VGND VGND VPWR VPWR _24149_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12094_ _12094_/A VGND VGND VPWR VPWR _12094_/Y sky130_fd_sc_hd__inv_2
X_16971_ _16021_/Y _24403_/Q _16021_/Y _24403_/Q VGND VGND VPWR VPWR _16972_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18710_ _18710_/A _18713_/A VGND VGND VPWR VPWR _18710_/X sky130_fd_sc_hd__and2_4
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15881__B1 _11766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15922_ _15922_/A VGND VGND VPWR VPWR _15923_/B sky130_fd_sc_hd__inv_2
X_19690_ _19688_/Y _19689_/X _19566_/X _19689_/X VGND VGND VPWR VPWR _23663_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18641_ _16627_/A _24133_/Q _16627_/Y _18689_/B VGND VGND VPWR VPWR _18641_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21905__A _21267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15853_ _15655_/X _15774_/X _15851_/X _21024_/B _15852_/X VGND VGND VPWR VPWR _15853_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_209_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15633__B1 _15632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14804_ _23983_/Q VGND VGND VPWR VPWR _14804_/Y sky130_fd_sc_hd__inv_2
X_18572_ _18476_/A _18572_/B VGND VGND VPWR VPWR _18573_/B sky130_fd_sc_hd__or2_4
X_12996_ _25361_/Q VGND VGND VPWR VPWR _12996_/Y sky130_fd_sc_hd__inv_2
X_15784_ _15560_/X _15659_/B VGND VGND VPWR VPWR _15784_/X sky130_fd_sc_hd__or2_4
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17523_ _25532_/Q _24303_/Q _11840_/Y _17522_/Y VGND VGND VPWR VPWR _17524_/D sky130_fd_sc_hd__o22a_4
XFILLER_91_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11947_ _19636_/A VGND VGND VPWR VPWR _11947_/Y sky130_fd_sc_hd__inv_2
X_14735_ _14734_/Y _14717_/X _14734_/A _14715_/X VGND VGND VPWR VPWR _14735_/X sky130_fd_sc_hd__o22a_4
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13423__A _13423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14666_ _14665_/Y VGND VGND VPWR VPWR _19054_/A sky130_fd_sc_hd__buf_2
X_17454_ _11656_/A _11660_/A _11979_/B VGND VGND VPWR VPWR _17484_/A sky130_fd_sc_hd__or3_4
X_11878_ _25523_/Q _11900_/A VGND VGND VPWR VPWR _11897_/A sky130_fd_sc_hd__and2_4
XFILLER_177_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13617_ _13635_/B VGND VGND VPWR VPWR _13617_/Y sky130_fd_sc_hd__inv_2
X_16405_ _24608_/Q VGND VGND VPWR VPWR _16405_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14597_ _14582_/A _14595_/X _14596_/X _13779_/X _25099_/Q VGND VGND VPWR VPWR _14597_/X
+ sky130_fd_sc_hd__a32o_4
X_17385_ _17391_/A _17391_/B VGND VGND VPWR VPWR _17389_/B sky130_fd_sc_hd__or2_4
XFILLER_220_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16734__A _16464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19124_ _19123_/Y _19121_/X _19008_/X _19121_/X VGND VGND VPWR VPWR _23859_/D sky130_fd_sc_hd__a2bb2o_4
X_13548_ _13548_/A VGND VGND VPWR VPWR _15701_/A sky130_fd_sc_hd__inv_2
X_16336_ _24632_/Q VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _16266_/Y _16264_/X _16073_/X _16264_/X VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__a2bb2o_4
X_19055_ _19054_/X VGND VGND VPWR VPWR _19061_/A sky130_fd_sc_hd__buf_2
XFILLER_185_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13479_ _13484_/C _13484_/D _13542_/C _12068_/X VGND VGND VPWR VPWR _13480_/A sky130_fd_sc_hd__or4_4
XFILLER_146_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15218_ _15251_/A _15248_/A _15073_/X _15172_/X VGND VGND VPWR VPWR _15218_/X sky130_fd_sc_hd__or4_4
X_18006_ _18006_/A VGND VGND VPWR VPWR _18090_/A sky130_fd_sc_hd__buf_2
X_16198_ _16189_/Y _16197_/X _11752_/X _16197_/X VGND VGND VPWR VPWR _16198_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15149_ _15370_/A _24600_/Q _15370_/A _24600_/Q VGND VGND VPWR VPWR _15150_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17565__A _17691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24088__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19957_ _19957_/A VGND VGND VPWR VPWR _21676_/B sky130_fd_sc_hd__inv_2
XANTENNA__24040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_222_0_HCLK clkbuf_8_222_0_HCLK/A VGND VGND VPWR VPWR _24602_/CLK sky130_fd_sc_hd__clkbuf_1
X_18908_ _14479_/A VGND VGND VPWR VPWR _18908_/X sky130_fd_sc_hd__buf_2
XANTENNA__19780__A _19765_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19888_ _19895_/A VGND VGND VPWR VPWR _19888_/X sky130_fd_sc_hd__buf_2
XANTENNA__12686__B1 _12662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12321__A2_N _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18839_ _16492_/Y _24153_/Q _16492_/Y _24153_/Q VGND VGND VPWR VPWR _18840_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21815__A _21815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15624__B1 _11834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21850_ _20525_/B _14203_/X _14275_/Y _21726_/B VGND VGND VPWR VPWR _21850_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20801_ _13145_/B _13144_/X VGND VGND VPWR VPWR _20801_/Y sky130_fd_sc_hd__nor2_4
X_21781_ _22390_/A _21781_/B _21780_/X VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__and3_4
XFILLER_36_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23520_ _25491_/CLK _20091_/X VGND VGND VPWR VPWR _13357_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20732_ _20730_/A _20725_/X _20731_/X VGND VGND VPWR VPWR _20732_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23451_ _24684_/CLK _23451_/D VGND VGND VPWR VPWR _23451_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20663_ _20663_/A VGND VGND VPWR VPWR _20663_/Y sky130_fd_sc_hd__inv_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22402_ _22014_/X VGND VGND VPWR VPWR _22402_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19020__A _19020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23382_ _21025_/X VGND VGND VPWR VPWR IRQ[26] sky130_fd_sc_hd__buf_2
XFILLER_137_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20594_ _14432_/Y _20574_/X _20564_/X _20593_/X VGND VGND VPWR VPWR _20594_/X sky130_fd_sc_hd__a211o_4
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24881__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25121_ _25154_/CLK _14498_/X HRESETn VGND VGND VPWR VPWR _25121_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22333_ _22333_/A VGND VGND VPWR VPWR _22333_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24810__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25052_ _24340_/CLK _14866_/X HRESETn VGND VGND VPWR VPWR _25052_/Q sky130_fd_sc_hd__dfrtp_4
X_22264_ _22264_/A _22264_/B VGND VGND VPWR VPWR _22265_/C sky130_fd_sc_hd__or2_4
XFILLER_133_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24003_ _24003_/CLK sda_i_S5 HRESETn VGND VGND VPWR VPWR _24004_/D sky130_fd_sc_hd__dfrtp_4
X_21215_ _21180_/X _21198_/X _21214_/X VGND VGND VPWR VPWR _21225_/B sky130_fd_sc_hd__and3_4
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22195_ _20518_/A _22176_/B _23980_/Q _21369_/B VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21709__B _23016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21146_ _12184_/A _12102_/X _12055_/Y _12102_/X VGND VGND VPWR VPWR _21146_/X sky130_fd_sc_hd__a2bb2o_4
X_21077_ _21058_/A _21069_/X _21077_/C VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__and3_4
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20028_ _23543_/Q VGND VGND VPWR VPWR _20028_/Y sky130_fd_sc_hd__inv_2
X_24905_ _24488_/CLK _15630_/X HRESETn VGND VGND VPWR VPWR _24905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_219_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15615__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _12850_/A _12780_/Y VGND VGND VPWR VPWR _12862_/C sky130_fd_sc_hd__or2_4
XANTENNA__15723__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24836_ _24825_/CLK _15834_/X HRESETn VGND VGND VPWR VPWR _24836_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21444__B _23016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11799_/Y _11794_/X _11800_/X _11794_/X VGND VGND VPWR VPWR _25542_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _24814_/Q VGND VGND VPWR VPWR _12781_/Y sky130_fd_sc_hd__inv_2
X_24767_ _24767_/CLK _15979_/X HRESETn VGND VGND VPWR VPWR _24767_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _14635_/Y _19610_/X _14622_/Y _19614_/A VGND VGND VPWR VPWR _21979_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14519_/X VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _12073_/A VGND VGND VPWR VPWR _11733_/B sky130_fd_sc_hd__inv_2
X_23718_ _23678_/CLK _19523_/X VGND VGND VPWR VPWR _19522_/A sky130_fd_sc_hd__dfxtp_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24698_ _24756_/CLK _16146_/X HRESETn VGND VGND VPWR VPWR _22649_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14446_/A VGND VGND VPWR VPWR _14451_/X sky130_fd_sc_hd__buf_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11663_/A _11663_/B _11663_/C VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__and3_4
X_23649_ _23644_/CLK _19729_/X VGND VGND VPWR VPWR _13333_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13217_/X _13400_/X _13402_/C VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__and3_4
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _17136_/X VGND VGND VPWR VPWR _17170_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _20477_/A VGND VGND VPWR VPWR _14382_/Y sky130_fd_sc_hd__inv_2
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16120_/Y _16116_/X _15960_/X _16116_/X VGND VGND VPWR VPWR _24708_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_229_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13333_ _13428_/A _13333_/B VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__or2_4
X_25319_ _25316_/CLK _13511_/X HRESETn VGND VGND VPWR VPWR _25319_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24551__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _16051_/Y _16049_/X _11818_/X _16049_/X VGND VGND VPWR VPWR _24734_/D sky130_fd_sc_hd__a2bb2o_4
X_13264_ _13171_/X _13259_/X _13264_/C VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__or3_4
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22291__A _24623_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15003_ _15003_/A VGND VGND VPWR VPWR _15182_/B sky130_fd_sc_hd__buf_2
X_12215_ _25462_/Q VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__inv_2
XANTENNA__17385__A _17391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13195_ _13195_/A _20422_/A VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__or2_4
XANTENNA__14802__A _14801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19811_ _19809_/Y _19806_/X _19810_/X _19806_/X VGND VGND VPWR VPWR _23622_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12146_ _12136_/B VGND VGND VPWR VPWR _12146_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19742_ _19741_/X VGND VGND VPWR VPWR _19742_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19045__B1 _18975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12077_ _12077_/A VGND VGND VPWR VPWR _21031_/A sky130_fd_sc_hd__buf_2
X_16954_ _16947_/X _16954_/B _16954_/C _16954_/D VGND VGND VPWR VPWR _16961_/C sky130_fd_sc_hd__or4_4
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21927__B1 _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15905_ _11830_/X VGND VGND VPWR VPWR _15905_/X sky130_fd_sc_hd__buf_2
XFILLER_110_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19673_ _13158_/B VGND VGND VPWR VPWR _19673_/Y sky130_fd_sc_hd__inv_2
X_16885_ _19800_/A VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__buf_2
XFILLER_38_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18624_ _24149_/Q VGND VGND VPWR VPWR _18765_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_52_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _24383_/CLK sky130_fd_sc_hd__clkbuf_1
X_15836_ _12314_/Y _15835_/X _11831_/X _15835_/X VGND VGND VPWR VPWR _15836_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18555_ _18554_/X VGND VGND VPWR VPWR _24177_/D sky130_fd_sc_hd__inv_2
X_12979_ _12853_/Y _12988_/B VGND VGND VPWR VPWR _12986_/B sky130_fd_sc_hd__or2_4
X_15767_ HWDATA[8] VGND VGND VPWR VPWR _15767_/X sky130_fd_sc_hd__buf_2
X_17506_ _11772_/Y _17572_/A _11772_/Y _17572_/A VGND VGND VPWR VPWR _17506_/X sky130_fd_sc_hd__a2bb2o_4
X_14718_ _14730_/C _14712_/X _14717_/X VGND VGND VPWR VPWR _14718_/Y sky130_fd_sc_hd__a21oi_4
X_18486_ _18516_/A _18486_/B _18486_/C _18486_/D VGND VGND VPWR VPWR _18486_/X sky130_fd_sc_hd__or4_4
XANTENNA__15071__C _15292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15698_ _15698_/A VGND VGND VPWR VPWR _15698_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17437_ _17436_/Y _17434_/X _16791_/X _17434_/X VGND VGND VPWR VPWR _24335_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14649_ _18051_/A VGND VGND VPWR VPWR _18016_/A sky130_fd_sc_hd__buf_2
XANTENNA__12992__A _24786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16464__A _16464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__B1 _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24639__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _17370_/B VGND VGND VPWR VPWR _17369_/B sky130_fd_sc_hd__inv_2
XFILLER_186_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19107_ _23865_/Q VGND VGND VPWR VPWR _21906_/B sky130_fd_sc_hd__inv_2
X_16319_ _24638_/Q VGND VGND VPWR VPWR _16319_/Y sky130_fd_sc_hd__inv_2
X_17299_ _17298_/X VGND VGND VPWR VPWR _17299_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19038_ _19036_/Y _19030_/X _19012_/X _19037_/X VGND VGND VPWR VPWR _19038_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_217_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_19_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21000_ _21000_/A _21000_/B VGND VGND VPWR VPWR _21000_/Y sky130_fd_sc_hd__nor2_4
XFILLER_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15845__B1 _24829_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22951_ _23020_/A _22938_/Y _22944_/X _22951_/D VGND VGND VPWR VPWR _22951_/X sky130_fd_sc_hd__or4_4
XFILLER_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21902_ _21897_/X _21901_/X _22214_/A VGND VGND VPWR VPWR _21902_/X sky130_fd_sc_hd__o21a_4
XFILLER_244_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20208__A2_N _20205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22882_ _22155_/B VGND VGND VPWR VPWR _22882_/X sky130_fd_sc_hd__buf_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16270__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24621_ _24625_/CLK _24621_/D HRESETn VGND VGND VPWR VPWR _21870_/A sky130_fd_sc_hd__dfrtp_4
X_21833_ _21817_/X _21832_/X _21511_/X VGND VGND VPWR VPWR _21833_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24552_ _24552_/CLK _24552_/D HRESETn VGND VGND VPWR VPWR _24552_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21764_ _21783_/A _19268_/Y VGND VGND VPWR VPWR _21764_/X sky130_fd_sc_hd__or2_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22894__B2 _21229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16022__B1 _11773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23503_ _23926_/CLK _23503_/D VGND VGND VPWR VPWR _20140_/A sky130_fd_sc_hd__dfxtp_4
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20715_ _20715_/A VGND VGND VPWR VPWR _20715_/Y sky130_fd_sc_hd__inv_2
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24483_ _24981_/CLK _16735_/X HRESETn VGND VGND VPWR VPWR _24483_/Q sky130_fd_sc_hd__dfrtp_4
X_21695_ _21468_/X _21695_/B VGND VGND VPWR VPWR _21696_/C sky130_fd_sc_hd__or2_4
XFILLER_51_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16374__A _24617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23434_ _23555_/CLK _23434_/D VGND VGND VPWR VPWR _20326_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20646_ _20622_/Y VGND VGND VPWR VPWR _20646_/X sky130_fd_sc_hd__buf_2
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23365_ VGND VGND VPWR VPWR _23365_/HI IRQ[29] sky130_fd_sc_hd__conb_1
XANTENNA__15128__A2 _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20577_ _14441_/Y _20574_/X _20565_/X _20576_/X VGND VGND VPWR VPWR _20578_/A sky130_fd_sc_hd__a211o_4
XFILLER_192_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25104_ _25105_/CLK _14559_/X HRESETn VGND VGND VPWR VPWR _25104_/Q sky130_fd_sc_hd__dfrtp_4
X_22316_ _15114_/A _22316_/B VGND VGND VPWR VPWR _22319_/B sky130_fd_sc_hd__or2_4
X_23296_ _23296_/A _23296_/B VGND VGND VPWR VPWR _23296_/X sky130_fd_sc_hd__or2_4
XANTENNA__14887__A1 _14885_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12843__A2_N _22302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25035_ _25030_/CLK _25035_/D HRESETn VGND VGND VPWR VPWR _25035_/Q sky130_fd_sc_hd__dfrtp_4
X_22247_ _22260_/A _22247_/B VGND VGND VPWR VPWR _22247_/X sky130_fd_sc_hd__or2_4
XFILLER_117_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15718__A _15718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15140__A2_N _16427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ _20971_/A _12000_/B VGND VGND VPWR VPWR _12000_/X sky130_fd_sc_hd__and2_4
XANTENNA__16089__B1 _24719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22178_ _22177_/X VGND VGND VPWR VPWR _22178_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15836__B1 _11831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21129_ _11744_/X VGND VGND VPWR VPWR _21129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13238__A _13322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21455__A _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13951_ _13951_/A _13951_/B _13935_/X _13967_/C VGND VGND VPWR VPWR _13952_/D sky130_fd_sc_hd__or4_4
XANTENNA__20963__A1_N _20836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ _12780_/Y _12906_/B _12883_/X _12899_/B VGND VGND VPWR VPWR _12902_/X sky130_fd_sc_hd__a211o_4
XFILLER_19_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13882_ _13880_/X _13881_/X _14272_/A _13876_/X VGND VGND VPWR VPWR _13882_/X sky130_fd_sc_hd__o22a_4
X_16670_ _16669_/Y _16667_/X _16402_/X _16667_/X VGND VGND VPWR VPWR _16670_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12833_ _24812_/Q VGND VGND VPWR VPWR _12833_/Y sky130_fd_sc_hd__inv_2
X_15621_ _15626_/A VGND VGND VPWR VPWR _15621_/X sky130_fd_sc_hd__buf_2
X_24819_ _24803_/CLK _24819_/D HRESETn VGND VGND VPWR VPWR _24819_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18340_ _20079_/C _17497_/Y _19075_/B _18333_/B VGND VGND VPWR VPWR _24214_/D sky130_fd_sc_hd__o22a_4
X_12764_ _22564_/A VGND VGND VPWR VPWR _12764_/Y sky130_fd_sc_hd__inv_2
X_15552_ _15551_/Y _15547_/X HADDR[0] _15547_/X VGND VGND VPWR VPWR _24930_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_199_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16013__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22286__A _22425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _25556_/Q VGND VGND VPWR VPWR _11715_/Y sky130_fd_sc_hd__inv_2
X_14503_ _13985_/X VGND VGND VPWR VPWR _14550_/A sky130_fd_sc_hd__buf_2
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _14412_/A VGND VGND VPWR VPWR _15483_/X sky130_fd_sc_hd__buf_2
X_18271_ _23358_/A _18270_/Y _16791_/X _18270_/Y VGND VGND VPWR VPWR _24230_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22717__C _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12695_ _12680_/A _12689_/B _12695_/C VGND VGND VPWR VPWR _12695_/X sky130_fd_sc_hd__and3_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16284__A _15681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24732__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _16314_/Y _17310_/A _16314_/Y _17310_/A VGND VGND VPWR VPWR _17222_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _25145_/Q VGND VGND VPWR VPWR _14434_/Y sky130_fd_sc_hd__inv_2
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _14354_/B VGND VGND VPWR VPWR _14365_/X sky130_fd_sc_hd__buf_2
X_17153_ _16987_/Y _17157_/A VGND VGND VPWR VPWR _17153_/Y sky130_fd_sc_hd__nand2_4
XFILLER_128_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13385_/A _13316_/B VGND VGND VPWR VPWR _13316_/X sky130_fd_sc_hd__or2_4
X_16104_ _16103_/X VGND VGND VPWR VPWR _16104_/X sky130_fd_sc_hd__buf_2
XFILLER_171_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17084_ _17393_/B _17080_/B _17083_/X VGND VGND VPWR VPWR _17084_/X sky130_fd_sc_hd__or3_4
XFILLER_155_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14296_ _14296_/A VGND VGND VPWR VPWR _14300_/A sky130_fd_sc_hd__inv_2
XFILLER_143_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13247_ _13242_/X _13244_/X _13246_/X VGND VGND VPWR VPWR _13247_/X sky130_fd_sc_hd__and3_4
X_16035_ _24740_/Q VGND VGND VPWR VPWR _16035_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ _13178_/A VGND VGND VPWR VPWR _13198_/A sky130_fd_sc_hd__buf_2
XANTENNA__20415__A3 _15993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13793__D _13793_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15827__B1 _24841_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12127_/Y _12123_/X _11867_/X _12128_/X VGND VGND VPWR VPWR _12129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19018__B1 _18991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17986_ _18008_/A VGND VGND VPWR VPWR _17987_/A sky130_fd_sc_hd__buf_2
XFILLER_229_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19725_ _19719_/Y VGND VGND VPWR VPWR _19725_/X sky130_fd_sc_hd__buf_2
X_16937_ _16937_/A VGND VGND VPWR VPWR _16937_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12987__A _21035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19656_ _19148_/A VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__buf_2
X_16868_ _14791_/X VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__buf_2
XANTENNA__15055__B2 _15024_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18607_ _16550_/Y _18606_/X _16550_/Y _24162_/Q VGND VGND VPWR VPWR _18612_/B sky130_fd_sc_hd__a2bb2o_4
X_15819_ _12317_/Y _15818_/X _11787_/X _15818_/X VGND VGND VPWR VPWR _15819_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_241_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19587_ _19574_/Y VGND VGND VPWR VPWR _19587_/X sky130_fd_sc_hd__buf_2
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16799_ _24452_/Q VGND VGND VPWR VPWR _16799_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21128__B2 _15674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18538_ _18471_/D _18538_/B VGND VGND VPWR VPWR _18539_/B sky130_fd_sc_hd__or2_4
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18469_ _24178_/Q VGND VGND VPWR VPWR _18539_/A sky130_fd_sc_hd__inv_2
XFILLER_221_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _20525_/A _15446_/A _20498_/X _15446_/A _20499_/X VGND VGND VPWR VPWR _20501_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_193_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21480_ _21474_/A _21480_/B VGND VGND VPWR VPWR _21480_/X sky130_fd_sc_hd__or2_4
XFILLER_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11919__A2 _11889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _20429_/Y _20430_/X _20243_/X _20430_/X VGND VGND VPWR VPWR _20431_/X sky130_fd_sc_hd__a2bb2o_4
X_23150_ _24545_/Q _22940_/X _22941_/X _23149_/X VGND VGND VPWR VPWR _23151_/C sky130_fd_sc_hd__a211o_4
X_20362_ _20362_/A VGND VGND VPWR VPWR _20362_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22101_ _21278_/X _22062_/Y _22067_/X _21519_/X _22100_/X VGND VGND VPWR VPWR _22101_/X
+ sky130_fd_sc_hd__a32o_4
X_23081_ _16754_/A _23016_/X _22903_/X VGND VGND VPWR VPWR _23081_/X sky130_fd_sc_hd__o21a_4
XFILLER_228_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15538__A _15544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20293_ _23446_/Q VGND VGND VPWR VPWR _21414_/B sky130_fd_sc_hd__inv_2
XANTENNA__14442__A _14442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22032_ _22032_/A _20021_/Y VGND VGND VPWR VPWR _22032_/X sky130_fd_sc_hd__or2_4
XFILLER_103_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12344__A2 _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19009__B1 _19008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16491__B1 _16315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20147__A2_N _20141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23983_ _24343_/CLK _23983_/D HRESETn VGND VGND VPWR VPWR _23983_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22934_ _22934_/A _23140_/B VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__and2_4
XFILLER_228_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16243__B1 _16241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21425__D _21425_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22865_ _16132_/Y _22531_/B _15870_/B _11799_/Y _22864_/X VGND VGND VPWR VPWR _22865_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_243_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13505__B _12107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21816_ _21812_/X _21815_/X _18306_/X VGND VGND VPWR VPWR _21817_/C sky130_fd_sc_hd__o21a_4
X_24604_ _24602_/CLK _24604_/D HRESETn VGND VGND VPWR VPWR _24604_/Q sky130_fd_sc_hd__dfrtp_4
X_22796_ _22436_/X _22781_/X _22786_/X _22795_/X VGND VGND VPWR VPWR _22796_/X sky130_fd_sc_hd__or4_4
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24535_ _24566_/CLK _24535_/D HRESETn VGND VGND VPWR VPWR _16594_/A sky130_fd_sc_hd__dfrtp_4
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21747_ _21747_/A VGND VGND VPWR VPWR _22941_/A sky130_fd_sc_hd__buf_2
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ _12218_/Y _12278_/Y _12238_/Y _12502_/A VGND VGND VPWR VPWR _12480_/X sky130_fd_sc_hd__or4_4
X_24466_ _24430_/CLK _24466_/D HRESETn VGND VGND VPWR VPWR _16770_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_200_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21678_ _21674_/X _21677_/X _18306_/X VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__o21a_4
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23684_/CLK _20371_/X VGND VGND VPWR VPWR _20369_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20629_ _17398_/B _20627_/Y _20628_/X VGND VGND VPWR VPWR _20629_/X sky130_fd_sc_hd__and3_4
XFILLER_184_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24397_ _24407_/CLK _17113_/X HRESETn VGND VGND VPWR VPWR _24397_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16453__A2_N _16384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14150_ _23967_/D _14149_/Y _25146_/Q _23967_/D VGND VGND VPWR VPWR _25226_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18750__C _18733_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23348_ _23188_/X _23345_/X _23347_/X VGND VGND VPWR VPWR _23348_/X sky130_fd_sc_hd__and3_4
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13101_ _12339_/Y _13104_/B VGND VGND VPWR VPWR _13102_/C sky130_fd_sc_hd__nand2_4
XFILLER_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11791__B1 _11790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14081_ _14045_/C _14543_/B VGND VGND VPWR VPWR _14082_/B sky130_fd_sc_hd__nor2_4
X_23279_ _12226_/Y _22444_/X _22730_/X _12337_/Y _22858_/X VGND VGND VPWR VPWR _23279_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__25349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13032_ _13026_/C _13029_/X VGND VGND VPWR VPWR _13032_/X sky130_fd_sc_hd__or2_4
X_25018_ _25018_/CLK _15283_/X HRESETn VGND VGND VPWR VPWR _15282_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_140_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15809__B1 _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17840_ _17766_/B _17818_/X VGND VGND VPWR VPWR _17843_/B sky130_fd_sc_hd__or2_4
XFILLER_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15094__A2_N _24601_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23347__A2 _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17771_ _17771_/A _16952_/Y _17753_/X _17770_/X VGND VGND VPWR VPWR _17771_/X sky130_fd_sc_hd__or4_4
X_14983_ _14983_/A _14983_/B _14983_/C _14982_/X VGND VGND VPWR VPWR _14983_/X sky130_fd_sc_hd__or4_4
XFILLER_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22555__B1 _22431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19510_ _23723_/Q VGND VGND VPWR VPWR _22267_/B sky130_fd_sc_hd__inv_2
XFILLER_219_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16722_ _16720_/Y _16716_/X _16368_/X _16721_/X VGND VGND VPWR VPWR _24487_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ _13934_/A VGND VGND VPWR VPWR _13934_/X sky130_fd_sc_hd__buf_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19441_ _17995_/B VGND VGND VPWR VPWR _19441_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21913__A _14709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16653_ _16653_/A VGND VGND VPWR VPWR _16709_/A sky130_fd_sc_hd__buf_2
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13865_ _24007_/Q VGND VGND VPWR VPWR _13876_/A sky130_fd_sc_hd__inv_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24913__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ _24915_/Q VGND VGND VPWR VPWR _15604_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12816_ _22678_/A _22669_/A _22678_/A _22669_/A VGND VGND VPWR VPWR _12824_/A sky130_fd_sc_hd__a2bb2o_4
X_19372_ _19371_/Y _19369_/X _19305_/X _19369_/X VGND VGND VPWR VPWR _19372_/X sky130_fd_sc_hd__a2bb2o_4
X_16584_ _16584_/A VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__buf_2
X_13796_ _11731_/A VGND VGND VPWR VPWR _21140_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_126_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _24437_/CLK sky130_fd_sc_hd__clkbuf_1
X_18323_ _18306_/A _18301_/B _18302_/Y VGND VGND VPWR VPWR _18323_/X sky130_fd_sc_hd__o21a_4
X_15535_ _11740_/A VGND VGND VPWR VPWR _15653_/A sky130_fd_sc_hd__inv_2
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12747_ _12538_/Y _12647_/D _12657_/A _12745_/B VGND VGND VPWR VPWR _12747_/X sky130_fd_sc_hd__a211o_4
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_189_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25223_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_187_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13431__A _13315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18254_ _22550_/A _18252_/X _11830_/X _18252_/X VGND VGND VPWR VPWR _24241_/D sky130_fd_sc_hd__a2bb2o_4
X_12678_ _25427_/Q _12678_/B VGND VGND VPWR VPWR _12680_/B sky130_fd_sc_hd__or2_4
X_15466_ _13927_/B _20620_/A _15440_/X _13923_/A _15461_/X VGND VGND VPWR VPWR _15466_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _24355_/Q VGND VGND VPWR VPWR _17205_/Y sky130_fd_sc_hd__inv_2
X_14417_ _14417_/A _14416_/X VGND VGND VPWR VPWR _14428_/A sky130_fd_sc_hd__nor2_4
X_18185_ _18084_/X _18996_/A VGND VGND VPWR VPWR _18186_/C sky130_fd_sc_hd__or2_4
XANTENNA__23283__A1 _21456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15397_ _15310_/A _15424_/A _15423_/A _15423_/B VGND VGND VPWR VPWR _15397_/X sky130_fd_sc_hd__or4_4
XANTENNA__16742__A _16737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17136_ _17032_/Y _17052_/Y VGND VGND VPWR VPWR _17136_/X sky130_fd_sc_hd__or2_4
X_14348_ _25167_/Q VGND VGND VPWR VPWR _14349_/C sky130_fd_sc_hd__inv_2
XFILLER_116_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16593__A1_N _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14279_ _25192_/Q VGND VGND VPWR VPWR _14279_/Y sky130_fd_sc_hd__inv_2
X_17067_ _17067_/A VGND VGND VPWR VPWR _24408_/D sky130_fd_sc_hd__inv_2
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16018_ _16018_/A VGND VGND VPWR VPWR _16018_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16473__B1 _16294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17969_ _18069_/A _17961_/X _17968_/X _15686_/X _15694_/X VGND VGND VPWR VPWR _17969_/X
+ sky130_fd_sc_hd__o32a_4
X_19708_ _13362_/B VGND VGND VPWR VPWR _19708_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19411__B1 _19410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20980_ _12147_/X _12168_/X VGND VGND VPWR VPWR _20980_/X sky130_fd_sc_hd__and2_4
XFILLER_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16225__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19639_ _19639_/A VGND VGND VPWR VPWR _19639_/X sky130_fd_sc_hd__buf_2
XFILLER_226_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21823__A _22029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_22_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24654__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_85_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22650_ _22562_/X _22649_/X _22144_/A _11820_/A _22940_/A VGND VGND VPWR VPWR _22650_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21601_ _21295_/A VGND VGND VPWR VPWR _22298_/A sky130_fd_sc_hd__buf_2
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22581_ _21063_/A _22576_/X _21844_/X _22580_/Y VGND VGND VPWR VPWR _22582_/A sky130_fd_sc_hd__a211o_4
XANTENNA__14437__A _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24320_ _24327_/CLK _17627_/X HRESETn VGND VGND VPWR VPWR _24320_/Q sky130_fd_sc_hd__dfrtp_4
X_21532_ _22202_/C VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__buf_2
XANTENNA__14539__B1 _25107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23985__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24251_ _24252_/CLK _24251_/D HRESETn VGND VGND VPWR VPWR _24251_/Q sky130_fd_sc_hd__dfrtp_4
X_21463_ _21463_/A VGND VGND VPWR VPWR _21679_/A sky130_fd_sc_hd__buf_2
XFILLER_193_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19478__B1 _19410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23202_ _24644_/Q _21536_/X VGND VGND VPWR VPWR _23202_/X sky130_fd_sc_hd__or2_4
X_20414_ _20413_/Y _20411_/Y _20243_/X _20411_/Y VGND VGND VPWR VPWR _23400_/D sky130_fd_sc_hd__a2bb2o_4
X_24182_ _24552_/CLK _24182_/D HRESETn VGND VGND VPWR VPWR _24182_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21394_ _21408_/A _21394_/B VGND VGND VPWR VPWR _21394_/X sky130_fd_sc_hd__or2_4
XFILLER_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23133_ _12428_/A _22998_/X _17752_/A _22924_/X VGND VGND VPWR VPWR _23133_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11796__A _25543_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20345_ _17458_/C _20344_/X VGND VGND VPWR VPWR _20345_/X sky130_fd_sc_hd__or2_4
XFILLER_161_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23064_ _22787_/X _23060_/Y _22881_/X _23063_/X VGND VGND VPWR VPWR _23064_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14711__B1 _14709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20276_ _20276_/A VGND VGND VPWR VPWR _22385_/B sky130_fd_sc_hd__inv_2
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22785__B1 _24876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22015_ _21996_/C _20344_/X VGND VGND VPWR VPWR _22015_/Y sky130_fd_sc_hd__nor2_4
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15740__A1_N _12595_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22537__B1 _22516_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18205__A1 _17973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11980_ _11978_/Y _11979_/X _11976_/X VGND VGND VPWR VPWR _11980_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_124_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23966_ _23946_/CLK _23966_/D HRESETn VGND VGND VPWR VPWR _23966_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16216__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22829__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22917_ _24636_/Q _23165_/B VGND VGND VPWR VPWR _22917_/X sky130_fd_sc_hd__or2_4
X_23897_ _23880_/CLK _23897_/D VGND VGND VPWR VPWR _23897_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_204_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21760__B2 _21607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _14299_/B _13532_/X _25306_/Q VGND VGND VPWR VPWR _13650_/X sky130_fd_sc_hd__o21a_4
X_22848_ _22848_/A VGND VGND VPWR VPWR _22848_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A VGND VGND VPWR VPWR _12601_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22304__A3 _22303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13581_ _25263_/Q VGND VGND VPWR VPWR _13581_/Y sky130_fd_sc_hd__inv_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14992__D _14991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22779_ _21316_/X VGND VGND VPWR VPWR _22779_/X sky130_fd_sc_hd__buf_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12532_ _24870_/Q VGND VGND VPWR VPWR _12532_/Y sky130_fd_sc_hd__inv_2
X_15320_ _15319_/X VGND VGND VPWR VPWR _15321_/B sky130_fd_sc_hd__inv_2
XFILLER_169_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24518_ _24684_/CLK _16642_/X HRESETn VGND VGND VPWR VPWR _24518_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25498_ _24171_/CLK _25498_/D HRESETn VGND VGND VPWR VPWR _25498_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17192__A1 _24635_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17192__B2 _17331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12463_ _12257_/A _12462_/Y VGND VGND VPWR VPWR _12463_/X sky130_fd_sc_hd__or2_4
X_15251_ _15251_/A _15249_/A VGND VGND VPWR VPWR _15252_/C sky130_fd_sc_hd__or2_4
XANTENNA__19469__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24449_ _25043_/CLK _16809_/X HRESETn VGND VGND VPWR VPWR _24449_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14202_ _21861_/A VGND VGND VPWR VPWR _14202_/X sky130_fd_sc_hd__buf_2
X_15182_ _15182_/A _15182_/B _15181_/X VGND VGND VPWR VPWR _15182_/X sky130_fd_sc_hd__or3_4
X_12394_ _12225_/Y _12401_/B _12275_/Y _12394_/D VGND VGND VPWR VPWR _12395_/A sky130_fd_sc_hd__or4_4
XFILLER_126_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11764__B1 _11763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14133_ _14133_/A VGND VGND VPWR VPWR _14153_/A sky130_fd_sc_hd__buf_2
X_19990_ _19990_/A VGND VGND VPWR VPWR _19990_/X sky130_fd_sc_hd__buf_2
XFILLER_126_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14064_ _14543_/A _13985_/X _14069_/A _14063_/Y VGND VGND VPWR VPWR _14064_/X sky130_fd_sc_hd__o22a_4
X_18941_ _18936_/Y _18940_/X _17427_/X _18940_/X VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13015_ _13044_/A _13015_/B _13014_/X VGND VGND VPWR VPWR _13015_/X sky130_fd_sc_hd__and3_4
XFILLER_239_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17393__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18620__A1_N _16578_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18872_ _18856_/X _18861_/X _18872_/C _18872_/D VGND VGND VPWR VPWR _18872_/X sky130_fd_sc_hd__or4_4
XFILLER_95_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16455__B1 _16375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17823_ _16909_/A _17823_/B VGND VGND VPWR VPWR _17823_/X sky130_fd_sc_hd__or2_4
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13426__A _13282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ _24274_/Q VGND VGND VPWR VPWR _17864_/A sky130_fd_sc_hd__inv_2
XFILLER_236_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14966_ _15079_/A _16822_/A _14965_/A _16822_/A VGND VGND VPWR VPWR _14966_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16705_ _16703_/Y _16704_/X _16349_/X _16704_/X VGND VGND VPWR VPWR _16705_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13917_ _13978_/B _13916_/Y VGND VGND VPWR VPWR _13917_/X sky130_fd_sc_hd__or2_4
X_17685_ _17687_/A _17678_/X _17685_/C VGND VGND VPWR VPWR _17685_/X sky130_fd_sc_hd__and3_4
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14897_ _14897_/A VGND VGND VPWR VPWR _15178_/A sky130_fd_sc_hd__inv_2
XANTENNA__16737__A _16468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19424_ _18080_/B VGND VGND VPWR VPWR _19424_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15641__A _15626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16636_ _13751_/Y _16182_/B _16643_/B VGND VGND VPWR VPWR _16636_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _13848_/A VGND VGND VPWR VPWR _13848_/X sky130_fd_sc_hd__buf_2
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16975__A2_N _17050_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19355_ _18093_/B VGND VGND VPWR VPWR _19355_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19272__A2_N _19271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16567_ _16584_/A VGND VGND VPWR VPWR _16567_/X sky130_fd_sc_hd__buf_2
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13779_ _14611_/A VGND VGND VPWR VPWR _13779_/X sky130_fd_sc_hd__buf_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18952__A _18952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18306_ _18306_/A VGND VGND VPWR VPWR _18306_/X sky130_fd_sc_hd__buf_2
XANTENNA__13161__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15518_ _15517_/Y _15513_/X HADDR[15] _15513_/X VGND VGND VPWR VPWR _24945_/D sky130_fd_sc_hd__a2bb2o_4
X_19286_ _19280_/Y VGND VGND VPWR VPWR _19286_/X sky130_fd_sc_hd__buf_2
X_16498_ _16497_/Y _16495_/X _16412_/X _16495_/X VGND VGND VPWR VPWR _24572_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22474__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18237_ _17973_/A _18236_/X _24247_/Q _18031_/A VGND VGND VPWR VPWR _24247_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17568__A _17567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15449_ _13942_/X _15446_/X _15441_/X _13933_/X _15447_/X VGND VGND VPWR VPWR _15449_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16930__A1 _21531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18168_ _18168_/A _18168_/B VGND VGND VPWR VPWR _18168_/X sky130_fd_sc_hd__or2_4
XFILLER_144_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17119_ _17106_/A _17119_/B _17119_/C VGND VGND VPWR VPWR _24395_/D sky130_fd_sc_hd__and3_4
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18099_ _18164_/A _23849_/Q VGND VGND VPWR VPWR _18101_/B sky130_fd_sc_hd__or2_4
X_20130_ _22382_/B _20129_/X _20102_/X _20129_/X VGND VGND VPWR VPWR _20130_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20061_ _20057_/Y _20060_/X _19790_/X _20060_/X VGND VGND VPWR VPWR _23532_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22519__B1 _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13336__A _13153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21990__B2 _21991_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24835__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23820_ _24214_/CLK _23820_/D VGND VGND VPWR VPWR _19232_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_239_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23751_ _23735_/CLK _23751_/D VGND VGND VPWR VPWR _18149_/B sky130_fd_sc_hd__dfxtp_4
X_20963_ _20836_/X _20962_/X _24513_/Q _20883_/A VGND VGND VPWR VPWR _24076_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_241_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22702_ _22443_/A VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__buf_2
XFILLER_242_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _23799_/CLK _23682_/D VGND VGND VPWR VPWR _23682_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _20878_/X _20893_/X _16696_/A _20883_/X VGND VGND VPWR VPWR _20894_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22633_ _13671_/A _21320_/A _13141_/A _21322_/X VGND VGND VPWR VPWR _22633_/Y sky130_fd_sc_hd__a22oi_4
X_25421_ _25425_/CLK _25421_/D HRESETn VGND VGND VPWR VPWR _25421_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25352_ _25365_/CLK _13087_/Y HRESETn VGND VGND VPWR VPWR _12356_/A sky130_fd_sc_hd__dfrtp_4
X_22564_ _22564_/A _21104_/B VGND VGND VPWR VPWR _22564_/X sky130_fd_sc_hd__or2_4
XFILLER_139_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_172_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23454_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21515_ _23421_/Q _20343_/X _23397_/Q _19597_/X VGND VGND VPWR VPWR _21515_/X sky130_fd_sc_hd__o22a_4
X_24303_ _24302_/CLK _17689_/X HRESETn VGND VGND VPWR VPWR _24303_/Q sky130_fd_sc_hd__dfrtp_4
X_25283_ _23516_/CLK _25283_/D HRESETn VGND VGND VPWR VPWR _13766_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22495_ _21311_/A VGND VGND VPWR VPWR _22789_/B sky130_fd_sc_hd__buf_2
XFILLER_182_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16382__A _16382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_29_0_HCLK clkbuf_7_14_0_HCLK/X VGND VGND VPWR VPWR _24697_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16921__B2 _16920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24234_ _24238_/CLK _24234_/D HRESETn VGND VGND VPWR VPWR _24234_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21446_ _21235_/X VGND VGND VPWR VPWR _22530_/B sky130_fd_sc_hd__buf_2
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24165_ _24194_/CLK _18598_/X HRESETn VGND VGND VPWR VPWR _24165_/Q sky130_fd_sc_hd__dfrtp_4
X_21377_ _21369_/Y _21377_/B _21374_/X _21377_/D VGND VGND VPWR VPWR _21378_/B sky130_fd_sc_hd__and4_4
X_23116_ _23113_/X _23114_/X _22872_/X _24850_/Q _23115_/X VGND VGND VPWR VPWR _23116_/X
+ sky130_fd_sc_hd__a32o_4
X_20328_ _23433_/Q VGND VGND VPWR VPWR _20328_/Y sky130_fd_sc_hd__inv_2
X_24096_ _24095_/CLK _20545_/X HRESETn VGND VGND VPWR VPWR _20613_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12752__A1_N _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13499__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19808__A2_N _19806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23047_ _23042_/Y _23046_/Y _22868_/X VGND VGND VPWR VPWR _23047_/X sky130_fd_sc_hd__o21a_4
X_20259_ _20255_/Y _20258_/X _19817_/X _20258_/X VGND VGND VPWR VPWR _23460_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18102__A _18102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16437__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16988__A1 _16065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24576__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14820_ _14835_/A VGND VGND VPWR VPWR _14820_/X sky130_fd_sc_hd__buf_2
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24998_ _24981_/CLK _24998_/D HRESETn VGND VGND VPWR VPWR _24998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _22056_/A VGND VGND VPWR VPWR _14751_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11963_ _19900_/A VGND VGND VPWR VPWR _11963_/Y sky130_fd_sc_hd__inv_2
X_23949_ _23960_/CLK _23949_/D HRESETn VGND VGND VPWR VPWR _20552_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13702_ _13702_/A _13702_/B _11705_/A _25300_/Q VGND VGND VPWR VPWR _13703_/A sky130_fd_sc_hd__and4_4
XFILLER_245_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17470_ _18333_/C _13198_/A _18333_/C _13198_/A VGND VGND VPWR VPWR _17470_/X sky130_fd_sc_hd__a2bb2o_4
X_11894_ _11890_/X _11893_/X _11879_/A _11881_/X VGND VGND VPWR VPWR _11894_/X sky130_fd_sc_hd__a211o_4
X_14682_ _19142_/B _13610_/X _19166_/B VGND VGND VPWR VPWR _25076_/D sky130_fd_sc_hd__o21a_4
XFILLER_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16421_ _24601_/Q VGND VGND VPWR VPWR _16421_/Y sky130_fd_sc_hd__inv_2
X_13633_ _13611_/A VGND VGND VPWR VPWR _14667_/A sky130_fd_sc_hd__inv_2
XANTENNA__15180__B _15172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ _19138_/Y _19134_/X _19139_/X _19134_/A VGND VGND VPWR VPWR _23853_/D sky130_fd_sc_hd__a2bb2o_4
X_16352_ _16352_/A VGND VGND VPWR VPWR _16352_/X sky130_fd_sc_hd__buf_2
X_13564_ _13564_/A VGND VGND VPWR VPWR _13564_/Y sky130_fd_sc_hd__inv_2
X_15303_ _15303_/A _15347_/A VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__or2_4
X_12515_ _13017_/B VGND VGND VPWR VPWR _13051_/A sky130_fd_sc_hd__buf_2
X_19071_ _19070_/Y _19068_/X _19048_/X _19068_/X VGND VGND VPWR VPWR _23878_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23238__A1 _22563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13495_ _25325_/Q VGND VGND VPWR VPWR _13495_/Y sky130_fd_sc_hd__inv_2
X_16283_ _15664_/X _16288_/B _16090_/X _24650_/Q _16282_/X VGND VGND VPWR VPWR _24650_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14805__A scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16912__B2 _21066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18022_ _18063_/A _18022_/B _18021_/X VGND VGND VPWR VPWR _18027_/B sky130_fd_sc_hd__and3_4
XFILLER_185_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12446_ _12458_/A _12444_/X _12445_/X VGND VGND VPWR VPWR _25459_/D sky130_fd_sc_hd__and3_4
X_15234_ _15252_/A _15228_/X _15234_/C VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__and3_4
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12377_ _24847_/Q VGND VGND VPWR VPWR _12377_/Y sky130_fd_sc_hd__inv_2
X_15165_ _15164_/Y _16387_/A _15164_/Y _16387_/A VGND VGND VPWR VPWR _15165_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22461__A2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16676__B1 _16407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14116_ _14116_/A _14116_/B _14115_/X VGND VGND VPWR VPWR _14117_/A sky130_fd_sc_hd__or3_4
X_15096_ _25007_/Q VGND VGND VPWR VPWR _15096_/Y sky130_fd_sc_hd__inv_2
X_19973_ _22034_/B _19967_/X _19632_/X _19972_/X VGND VGND VPWR VPWR _19973_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22749__B1 _22431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18924_ _23929_/Q VGND VGND VPWR VPWR _21909_/B sky130_fd_sc_hd__inv_2
XANTENNA__15636__A _14427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14047_ _14047_/A VGND VGND VPWR VPWR _14060_/C sky130_fd_sc_hd__inv_2
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20224__B2 _20219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18855_ _24569_/Q _18764_/A _16522_/Y _24141_/Q VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22764__A3 _22157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ _17752_/A _17805_/Y VGND VGND VPWR VPWR _17806_/X sky130_fd_sc_hd__or2_4
XFILLER_227_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17851__A _17762_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18786_ _18786_/A VGND VGND VPWR VPWR _18786_/Y sky130_fd_sc_hd__inv_2
X_15998_ _15797_/X _15895_/A _15933_/X _21091_/A _15940_/X VGND VGND VPWR VPWR _24753_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23174__B1 _24289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ _18319_/A VGND VGND VPWR VPWR _17738_/A sky130_fd_sc_hd__buf_2
XFILLER_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14949_ _14905_/X _14919_/X _14949_/C _14948_/X VGND VGND VPWR VPWR _14994_/A sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_20_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22921__B1 _25544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17668_ _17687_/A _17666_/X _17668_/C VGND VGND VPWR VPWR _24309_/D sky130_fd_sc_hd__and3_4
XFILLER_51_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19407_ _18175_/B VGND VGND VPWR VPWR _19407_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16600__B1 _16245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16619_ _16617_/Y _16618_/X _16534_/X _16618_/X VGND VGND VPWR VPWR _24526_/D sky130_fd_sc_hd__a2bb2o_4
X_17599_ _17691_/A VGND VGND VPWR VPWR _17895_/B sky130_fd_sc_hd__inv_2
XFILLER_211_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19338_ _19324_/Y VGND VGND VPWR VPWR _19338_/X sky130_fd_sc_hd__buf_2
XANTENNA__17298__A _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_245_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _24981_/CLK sky130_fd_sc_hd__clkbuf_1
X_19269_ _19268_/Y _19264_/X _16890_/X _19264_/X VGND VGND VPWR VPWR _23808_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16903__B2 _17752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21300_ _21597_/A VGND VGND VPWR VPWR _21300_/Y sky130_fd_sc_hd__inv_2
X_22280_ _21288_/X _22242_/X _21968_/X _22279_/X VGND VGND VPWR VPWR _22281_/A sky130_fd_sc_hd__o22a_4
XFILLER_176_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22932__A _16682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21231_ _21231_/A VGND VGND VPWR VPWR _21877_/B sky130_fd_sc_hd__buf_2
X_21162_ _21004_/A _14201_/A _21160_/Y _21161_/X VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20113_ _21925_/B _20109_/X _20112_/X _20109_/X VGND VGND VPWR VPWR _23513_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21093_ _24786_/Q _15662_/Y _21049_/X _21092_/X VGND VGND VPWR VPWR _21093_/X sky130_fd_sc_hd__a211o_4
XFILLER_113_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20044_ _20038_/Y VGND VGND VPWR VPWR _20044_/X sky130_fd_sc_hd__buf_2
X_24921_ _24923_/CLK _24921_/D HRESETn VGND VGND VPWR VPWR _24921_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17761__A _16920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24852_ _24878_/CLK _15812_/X HRESETn VGND VGND VPWR VPWR _24852_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17631__A2 _17610_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23803_ _23514_/CLK _19284_/X VGND VGND VPWR VPWR _19283_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _18366_/Y _21995_/B VGND VGND VPWR VPWR _21995_/X sky130_fd_sc_hd__and2_4
X_24783_ _24803_/CLK _24783_/D HRESETn VGND VGND VPWR VPWR _24783_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20946_ _20927_/X _20945_/X _16666_/A _20931_/X VGND VGND VPWR VPWR _20946_/X sky130_fd_sc_hd__a2bb2o_4
X_23734_ _23735_/CLK _19476_/X VGND VGND VPWR VPWR _18184_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _20876_/X VGND VGND VPWR VPWR _24056_/D sky130_fd_sc_hd__inv_2
X_23665_ _23654_/CLK _19685_/X VGND VGND VPWR VPWR _13325_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_241_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_55_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25404_ _24799_/CLK _12870_/X HRESETn VGND VGND VPWR VPWR _25404_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _22616_/A _22578_/B VGND VGND VPWR VPWR _22616_/X sky130_fd_sc_hd__and2_4
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23596_ _23684_/CLK _23596_/D VGND VGND VPWR VPWR _23596_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22140__A1 _21547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22140__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22547_ _14909_/A _22541_/X _22542_/X _22546_/X VGND VGND VPWR VPWR _22547_/X sky130_fd_sc_hd__a211o_4
X_25335_ _25488_/CLK _25335_/D HRESETn VGND VGND VPWR VPWR _25335_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12300_ _12191_/Y _12414_/A VGND VGND VPWR VPWR _12393_/A sky130_fd_sc_hd__or2_4
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13280_ _13387_/A _13278_/X _13280_/C VGND VGND VPWR VPWR _13284_/B sky130_fd_sc_hd__and3_4
X_22478_ _20730_/Y _21605_/X _15625_/Y _22460_/X VGND VGND VPWR VPWR _22479_/B sky130_fd_sc_hd__o22a_4
X_25266_ _25309_/CLK _13847_/X HRESETn VGND VGND VPWR VPWR _25266_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ _12228_/A _22483_/A _12229_/X _12230_/Y VGND VGND VPWR VPWR _12231_/X sky130_fd_sc_hd__o22a_4
X_21429_ _21535_/A VGND VGND VPWR VPWR _22430_/A sky130_fd_sc_hd__buf_2
X_24217_ _24217_/CLK _24217_/D HRESETn VGND VGND VPWR VPWR _24217_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25197_ _25200_/CLK _14269_/X HRESETn VGND VGND VPWR VPWR _25197_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16658__B1 _16389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12162_ _12162_/A VGND VGND VPWR VPWR _12162_/Y sky130_fd_sc_hd__inv_2
X_24148_ _24989_/CLK _24148_/D HRESETn VGND VGND VPWR VPWR _18768_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21458__A _15792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24757__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12093_ _12092_/Y _12088_/X _11862_/X _12088_/X VGND VGND VPWR VPWR _25487_/D sky130_fd_sc_hd__a2bb2o_4
X_16970_ _24727_/Q _16969_/Y _16016_/Y _17080_/A VGND VGND VPWR VPWR _16970_/X sky130_fd_sc_hd__a2bb2o_4
X_24079_ _25365_/CLK _24079_/D HRESETn VGND VGND VPWR VPWR _24079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21891__A2_N _21890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15921_ _14778_/X _15919_/Y _15922_/A VGND VGND VPWR VPWR _15921_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20206__B2 _20205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18640_ _24133_/Q VGND VGND VPWR VPWR _18689_/B sky130_fd_sc_hd__inv_2
XANTENNA__17671__A _17567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15852_ _15659_/B _15854_/B VGND VGND VPWR VPWR _15852_/X sky130_fd_sc_hd__or2_4
XFILLER_49_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14803_ _13643_/A _13610_/X _14802_/Y _25062_/Q _14631_/Y VGND VGND VPWR VPWR _25062_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16830__B1 HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18571_ _18476_/B _18570_/X VGND VGND VPWR VPWR _18572_/B sky130_fd_sc_hd__or2_4
X_15783_ _15758_/X _15774_/X _15782_/X _24860_/Q _15719_/X VGND VGND VPWR VPWR _24860_/D
+ sky130_fd_sc_hd__a32o_4
X_12995_ _12308_/Y _12329_/Y VGND VGND VPWR VPWR _12995_/X sky130_fd_sc_hd__or2_4
XFILLER_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17522_ _24303_/Q VGND VGND VPWR VPWR _17522_/Y sky130_fd_sc_hd__inv_2
X_14734_ _14734_/A VGND VGND VPWR VPWR _14734_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11946_ _20000_/A VGND VGND VPWR VPWR _19636_/A sky130_fd_sc_hd__buf_2
XFILLER_189_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17453_ _17447_/Y _17450_/Y _17452_/X _17450_/Y VGND VGND VPWR VPWR _17453_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14665_ _25079_/Q VGND VGND VPWR VPWR _14665_/Y sky130_fd_sc_hd__inv_2
X_11877_ _11873_/Y _11750_/X _11876_/X _11750_/X VGND VGND VPWR VPWR _25525_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16404_ _15111_/Y _16398_/X _16402_/X _16403_/X VGND VGND VPWR VPWR _16404_/X sky130_fd_sc_hd__a2bb2o_4
X_13616_ _14794_/A _13614_/B _13615_/Y VGND VGND VPWR VPWR _13635_/B sky130_fd_sc_hd__o21a_4
X_17384_ _17384_/A VGND VGND VPWR VPWR _24350_/D sky130_fd_sc_hd__inv_2
X_14596_ _25099_/Q _14580_/A VGND VGND VPWR VPWR _14596_/X sky130_fd_sc_hd__or2_4
XFILLER_198_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19123_ _13215_/B VGND VGND VPWR VPWR _19123_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16945__A1_N _16138_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16734__B _16464_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16335_ _16331_/Y _16333_/X _16334_/X _16333_/X VGND VGND VPWR VPWR _24633_/D sky130_fd_sc_hd__a2bb2o_4
X_13547_ _13547_/A VGND VGND VPWR VPWR _13547_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19054_ _19054_/A _19143_/B _19054_/C _19054_/D VGND VGND VPWR VPWR _19054_/X sky130_fd_sc_hd__and4_4
X_16266_ _22107_/A VGND VGND VPWR VPWR _16266_/Y sky130_fd_sc_hd__inv_2
X_13478_ _13504_/B VGND VGND VPWR VPWR _13484_/D sky130_fd_sc_hd__buf_2
Xclkbuf_8_12_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23560_/CLK sky130_fd_sc_hd__clkbuf_1
X_18005_ _18102_/A VGND VGND VPWR VPWR _18127_/A sky130_fd_sc_hd__buf_2
X_15217_ _15293_/A VGND VGND VPWR VPWR _15252_/A sky130_fd_sc_hd__buf_2
X_12429_ _12398_/A _12429_/B _12429_/C VGND VGND VPWR VPWR _12429_/X sky130_fd_sc_hd__and3_4
XANTENNA__22434__A2 _22427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_75_0_HCLK clkbuf_8_74_0_HCLK/A VGND VGND VPWR VPWR _24756_/CLK sky130_fd_sc_hd__clkbuf_1
X_16197_ _16196_/X VGND VGND VPWR VPWR _16197_/X sky130_fd_sc_hd__buf_2
XFILLER_154_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19835__B1 _19761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15148_ _15383_/A VGND VGND VPWR VPWR _15370_/A sky130_fd_sc_hd__inv_2
XFILLER_126_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21368__A _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ _15079_/A _15009_/X _15069_/X _15078_/X VGND VGND VPWR VPWR _15080_/B sky130_fd_sc_hd__or4_4
X_19956_ _19955_/Y _19951_/X _19639_/X _19951_/X VGND VGND VPWR VPWR _23568_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18907_ _20430_/A VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__buf_2
X_19887_ _19887_/A VGND VGND VPWR VPWR _22026_/B sky130_fd_sc_hd__inv_2
X_18838_ _16542_/Y _24134_/Q _16542_/Y _24134_/Q VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22199__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16821__B1 HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18769_ _18776_/A _18769_/B _18769_/C VGND VGND VPWR VPWR _24148_/D sky130_fd_sc_hd__and3_4
XFILLER_215_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20800_ _20799_/X VGND VGND VPWR VPWR _24038_/D sky130_fd_sc_hd__inv_2
XFILLER_209_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21780_ _22090_/A _21780_/B VGND VGND VPWR VPWR _21780_/X sky130_fd_sc_hd__or2_4
XANTENNA__17377__A1 _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18574__B1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20731_ _20730_/Y _20731_/B VGND VGND VPWR VPWR _20731_/X sky130_fd_sc_hd__and2_4
XFILLER_91_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22646__B _22610_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23450_ _23475_/CLK _23450_/D VGND VGND VPWR VPWR _23450_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20662_ _14244_/Y _20646_/X _20637_/A _20661_/X VGND VGND VPWR VPWR _20663_/A sky130_fd_sc_hd__a211o_4
XFILLER_149_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22122__A1 _12952_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22401_ _22401_/A _22319_/X _22401_/C _22401_/D VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__or4_4
X_23381_ _21024_/X VGND VGND VPWR VPWR IRQ[25] sky130_fd_sc_hd__buf_2
X_20593_ _18886_/B _20592_/Y _20597_/C VGND VGND VPWR VPWR _20593_/X sky130_fd_sc_hd__and3_4
X_22332_ _21577_/X _22330_/X _21583_/X _22331_/X VGND VGND VPWR VPWR _22333_/A sky130_fd_sc_hd__o22a_4
X_25120_ _25154_/CLK _14500_/X HRESETn VGND VGND VPWR VPWR _14499_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_192_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22662__A _24630_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25051_ _24000_/CLK _25051_/D HRESETn VGND VGND VPWR VPWR _14823_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22263_ _18300_/B _19969_/Y VGND VGND VPWR VPWR _22265_/B sky130_fd_sc_hd__or2_4
XFILLER_247_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17756__A _21066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18629__A1 _16571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16660__A _16654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24002_ _24340_/CLK _24002_/D HRESETn VGND VGND VPWR VPWR _24002_/Q sky130_fd_sc_hd__dfrtp_4
X_21214_ _21463_/A _21205_/X _21213_/X VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__or3_4
XFILLER_183_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22194_ _22193_/X VGND VGND VPWR VPWR _22194_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24850__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21145_ _18901_/Y _21134_/Y _21348_/A _21144_/X VGND VGND VPWR VPWR _21226_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12126__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21076_ _21047_/X _21074_/X _21882_/A _21075_/X VGND VGND VPWR VPWR _21077_/C sky130_fd_sc_hd__a211o_4
XFILLER_120_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20027_ _21811_/B _20022_/X _20003_/X _20022_/X VGND VGND VPWR VPWR _20027_/X sky130_fd_sc_hd__a2bb2o_4
X_24904_ _24488_/CLK _15633_/X HRESETn VGND VGND VPWR VPWR _15631_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17491__A _17485_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16812__B1 HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24835_ _24878_/CLK _15836_/X HRESETn VGND VGND VPWR VPWR _24835_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ HWDATA[17] VGND VGND VPWR VPWR _11800_/X sky130_fd_sc_hd__buf_2
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13524__A _14248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _25397_/Q VGND VGND VPWR VPWR _12780_/Y sky130_fd_sc_hd__inv_2
X_24766_ _24757_/CLK _24766_/D HRESETn VGND VGND VPWR VPWR _22665_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _21975_/X _21976_/X _21977_/X VGND VGND VPWR VPWR _21978_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22837__A _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21741__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11731_/A _11731_/B VGND VGND VPWR VPWR _13822_/A sky130_fd_sc_hd__or2_4
X_23717_ _23717_/CLK _23717_/D VGND VGND VPWR VPWR _23717_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _13659_/A _24067_/Q _20907_/B _13658_/X VGND VGND VPWR VPWR _20929_/X sky130_fd_sc_hd__or4_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24697_ _24697_/CLK _24697_/D HRESETn VGND VGND VPWR VPWR _22613_/A sky130_fd_sc_hd__dfrtp_4
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14450_/A VGND VGND VPWR VPWR _14450_/Y sky130_fd_sc_hd__inv_2
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__inv_2
X_23648_ _23642_/CLK _23648_/D VGND VGND VPWR VPWR _13368_/B sky130_fd_sc_hd__dfxtp_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24094__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13369_/A _13401_/B VGND VGND VPWR VPWR _13402_/C sky130_fd_sc_hd__or2_4
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _25159_/Q _14369_/A _14365_/X _12099_/A _14364_/A VGND VGND VPWR VPWR _25159_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _23514_/CLK _19929_/X VGND VGND VPWR VPWR _23579_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _24708_/Q VGND VGND VPWR VPWR _16120_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13423_/A VGND VGND VPWR VPWR _13332_/X sky130_fd_sc_hd__buf_2
X_25318_ _25188_/CLK _13513_/X HRESETn VGND VGND VPWR VPWR _25318_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16051_ _16051_/A VGND VGND VPWR VPWR _16051_/Y sky130_fd_sc_hd__inv_2
X_13263_ _13177_/A _13260_/X _13263_/C VGND VGND VPWR VPWR _13264_/C sky130_fd_sc_hd__and3_4
X_25249_ _24138_/CLK _13892_/X HRESETn VGND VGND VPWR VPWR _21160_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_170_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22416__A2 _21113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22291__B _22291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15002_ _15002_/A VGND VGND VPWR VPWR _15003_/A sky130_fd_sc_hd__inv_2
X_12214_ _25446_/Q _12213_/A _12212_/X _12213_/Y VGND VGND VPWR VPWR _12214_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21624__B1 _14721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13194_ _13190_/X _13193_/X _13171_/X VGND VGND VPWR VPWR _13194_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24591__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _12125_/A _24113_/Q _12125_/A _24113_/Q VGND VGND VPWR VPWR _12145_/X sky130_fd_sc_hd__a2bb2o_4
X_19810_ _19810_/A VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__buf_2
XFILLER_123_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12117__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _11731_/B VGND VGND VPWR VPWR _13798_/B sky130_fd_sc_hd__buf_2
X_16953_ _24708_/Q _16952_/Y _16125_/Y _16950_/A VGND VGND VPWR VPWR _16954_/D sky130_fd_sc_hd__a2bb2o_4
X_19741_ _17463_/X _20079_/B _18959_/A _18959_/B VGND VGND VPWR VPWR _19741_/X sky130_fd_sc_hd__or4_4
XFILLER_238_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15904_ _15875_/Y VGND VGND VPWR VPWR _15904_/X sky130_fd_sc_hd__buf_2
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19672_ _19671_/Y _19667_/X _19620_/X _19652_/Y VGND VGND VPWR VPWR _23669_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16884_ _19803_/A VGND VGND VPWR VPWR _16884_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18623_ _18613_/X _18616_/X _18623_/C _18622_/X VGND VGND VPWR VPWR _18623_/X sky130_fd_sc_hd__or4_4
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ _15806_/Y VGND VGND VPWR VPWR _15835_/X sky130_fd_sc_hd__buf_2
XFILLER_64_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13434__A _13217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18554_ _18471_/D _18538_/B _18505_/X _18552_/B VGND VGND VPWR VPWR _18554_/X sky130_fd_sc_hd__a211o_4
X_15766_ _12558_/Y _15763_/X _15765_/X _15763_/X VGND VGND VPWR VPWR _24869_/D sky130_fd_sc_hd__a2bb2o_4
X_12978_ _12978_/A VGND VGND VPWR VPWR _25377_/D sky130_fd_sc_hd__inv_2
X_17505_ _25531_/Q _17504_/Y _11765_/Y _17512_/A VGND VGND VPWR VPWR _17507_/C sky130_fd_sc_hd__a2bb2o_4
X_14717_ _14716_/Y VGND VGND VPWR VPWR _14717_/X sky130_fd_sc_hd__buf_2
XANTENNA__21651__A _14725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11929_ _11929_/A VGND VGND VPWR VPWR _11929_/Y sky130_fd_sc_hd__inv_2
X_18485_ _18473_/X _18515_/B VGND VGND VPWR VPWR _18486_/D sky130_fd_sc_hd__or2_4
X_15697_ _15686_/X _15693_/A _14629_/B _15691_/C _15696_/X VGND VGND VPWR VPWR _15698_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12840__B2 _23290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17436_ _24335_/Q VGND VGND VPWR VPWR _17436_/Y sky130_fd_sc_hd__inv_2
X_14648_ _14794_/A VGND VGND VPWR VPWR _18051_/A sky130_fd_sc_hd__buf_2
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22104__A1 _14954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23301__B1 _25403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16464__B _16464_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11889__A _11889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _17364_/B _17364_/C VGND VGND VPWR VPWR _17370_/B sky130_fd_sc_hd__or2_4
X_14579_ _25098_/Q _14578_/Y VGND VGND VPWR VPWR _14580_/A sky130_fd_sc_hd__and2_4
XANTENNA__14265__A _21375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19106_ _22078_/B _19100_/X _16881_/X _19105_/X VGND VGND VPWR VPWR _23866_/D sky130_fd_sc_hd__a2bb2o_4
X_16318_ _16317_/Y _16312_/X _15960_/X _16312_/X VGND VGND VPWR VPWR _16318_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17298_ _17298_/A _17292_/Y _17297_/X VGND VGND VPWR VPWR _17298_/X sky130_fd_sc_hd__or3_4
X_19037_ _19037_/A VGND VGND VPWR VPWR _19037_/X sky130_fd_sc_hd__buf_2
XANTENNA__24679__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16249_ _16247_/Y _16242_/X _16248_/X _16242_/X VGND VGND VPWR VPWR _24664_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16480__A _24579_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24608__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14712__B _14713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15845__A1 _15833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15845__B2 _15802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19939_ _19937_/Y _19938_/X _19807_/X _19938_/X VGND VGND VPWR VPWR _23575_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13856__B1 _13524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22950_ _22950_/A _22946_/X _22950_/C VGND VGND VPWR VPWR _22951_/D sky130_fd_sc_hd__and3_4
XFILLER_56_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21901_ _22235_/A _21899_/X _21900_/X VGND VGND VPWR VPWR _21901_/X sky130_fd_sc_hd__and3_4
XFILLER_228_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22881_ _22204_/A VGND VGND VPWR VPWR _22881_/X sky130_fd_sc_hd__buf_2
XFILLER_244_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24620_ _24625_/CLK _16369_/X HRESETn VGND VGND VPWR VPWR _24620_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_241_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21832_ _22274_/A _21832_/B _21831_/X VGND VGND VPWR VPWR _21832_/X sky130_fd_sc_hd__or3_4
XANTENNA__14281__B1 _13812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21763_ _21644_/A _21763_/B VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__or2_4
X_24551_ _24562_/CLK _24551_/D HRESETn VGND VGND VPWR VPWR _16550_/A sky130_fd_sc_hd__dfrtp_4
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16655__A _16654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _15638_/Y _20695_/X _20704_/X _20713_/Y VGND VGND VPWR VPWR _20715_/A sky130_fd_sc_hd__o22a_4
X_23502_ _23926_/CLK _23502_/D VGND VGND VPWR VPWR _23502_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19031__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21694_ _21668_/A _21694_/B VGND VGND VPWR VPWR _21694_/X sky130_fd_sc_hd__or2_4
X_24482_ _25030_/CLK _16740_/X HRESETn VGND VGND VPWR VPWR _24482_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20645_ _20644_/X VGND VGND VPWR VPWR _23991_/D sky130_fd_sc_hd__inv_2
X_23433_ _23441_/CLK _23433_/D VGND VGND VPWR VPWR _23433_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23364_ VGND VGND VPWR VPWR _23364_/HI IRQ[28] sky130_fd_sc_hd__conb_1
X_20576_ _18881_/X _20575_/Y _20556_/X VGND VGND VPWR VPWR _20576_/X sky130_fd_sc_hd__and3_4
XFILLER_165_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25103_ _25103_/CLK _14585_/X HRESETn VGND VGND VPWR VPWR _25103_/Q sky130_fd_sc_hd__dfrtp_4
X_22315_ _16460_/A _22312_/X _22315_/C VGND VGND VPWR VPWR _22401_/A sky130_fd_sc_hd__and3_4
XFILLER_137_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17486__A _17485_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23295_ _23295_/A VGND VGND VPWR VPWR _23295_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16390__A _16390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20624__B _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22246_ _21685_/X _22244_/X _22245_/X VGND VGND VPWR VPWR _22246_/X sky130_fd_sc_hd__and3_4
X_25034_ _25030_/CLK _25034_/D HRESETn VGND VGND VPWR VPWR _15074_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22177_ _14448_/Y _14443_/A _14465_/Y _21373_/A VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21128_ _21048_/X _21127_/X _13150_/Y _15674_/A VGND VGND VPWR VPWR _21128_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13847__B1 _13846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15734__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13950_ _13950_/A VGND VGND VPWR VPWR _13950_/Y sky130_fd_sc_hd__inv_2
X_21059_ _24860_/Q _21039_/X _21042_/X _21058_/X VGND VGND VPWR VPWR _21060_/C sky130_fd_sc_hd__a211o_4
XFILLER_101_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12901_ _12906_/A _12901_/B _12901_/C VGND VGND VPWR VPWR _25398_/D sky130_fd_sc_hd__and3_4
XFILLER_235_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13881_ _22129_/A _13870_/X _21847_/A _13872_/X VGND VGND VPWR VPWR _13881_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12382__A2_N _24828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15620_ _24908_/Q VGND VGND VPWR VPWR _22577_/A sky130_fd_sc_hd__inv_2
XANTENNA__13254__A _13451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12832_ _12765_/Y _23162_/A _25393_/Q _12831_/Y VGND VGND VPWR VPWR _12836_/C sky130_fd_sc_hd__a2bb2o_4
X_24818_ _24803_/CLK _24818_/D HRESETn VGND VGND VPWR VPWR _23231_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15551_ _13603_/B VGND VGND VPWR VPWR _15551_/Y sky130_fd_sc_hd__inv_2
X_12763_ _12921_/C _24806_/Q _12921_/C _24806_/Q VGND VGND VPWR VPWR _12772_/A sky130_fd_sc_hd__a2bb2o_4
X_24749_ _24642_/CLK _24749_/D HRESETn VGND VGND VPWR VPWR _24749_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14501_/Y _14497_/X _14409_/X _14485_/A VGND VGND VPWR VPWR _25119_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_230_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11970_/C _11661_/X _11979_/B _11713_/Y VGND VGND VPWR VPWR _25557_/D sky130_fd_sc_hd__o22a_4
X_18270_ _18269_/X VGND VGND VPWR VPWR _18270_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _24959_/Q VGND VGND VPWR VPWR _15482_/Y sky130_fd_sc_hd__inv_2
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12618_/B _12685_/D VGND VGND VPWR VPWR _12695_/C sky130_fd_sc_hd__nand2_4
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_25_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _16341_/Y _17348_/A _16341_/Y _17348_/A VGND VGND VPWR VPWR _17225_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14432_/Y _14428_/X _14412_/X _14428_/X VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _17127_/X _17142_/X _17152_/C VGND VGND VPWR VPWR _17152_/X sky130_fd_sc_hd__and3_4
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _14364_/A VGND VGND VPWR VPWR _14364_/X sky130_fd_sc_hd__buf_2
XFILLER_11_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19595__B _21161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _16096_/X VGND VGND VPWR VPWR _16103_/X sky130_fd_sc_hd__buf_2
XANTENNA__24772__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _13315_/A _13315_/B _13314_/X VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__or3_4
X_17083_ _17057_/X _17074_/X _17035_/Y VGND VGND VPWR VPWR _17083_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14295_ _25188_/Q _14310_/A VGND VGND VPWR VPWR _25188_/D sky130_fd_sc_hd__and2_4
XFILLER_182_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24701__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16034_ _16033_/Y _16031_/X _15965_/X _16031_/X VGND VGND VPWR VPWR _24741_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13246_ _13245_/X _23659_/Q VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__or2_4
XFILLER_170_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13177_ _13177_/A VGND VGND VPWR VPWR _13200_/A sky130_fd_sc_hd__buf_2
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12333__A _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_149_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _24354_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12128_ _12123_/A VGND VGND VPWR VPWR _12128_/X sky130_fd_sc_hd__buf_2
X_17985_ _17985_/A VGND VGND VPWR VPWR _18008_/A sky130_fd_sc_hd__buf_2
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12059_ _12059_/A VGND VGND VPWR VPWR _16378_/A sky130_fd_sc_hd__buf_2
X_16936_ _17759_/C VGND VGND VPWR VPWR _16936_/X sky130_fd_sc_hd__buf_2
X_19724_ _13295_/B VGND VGND VPWR VPWR _19724_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18020__A _18013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12987__B _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16867_ _16866_/X VGND VGND VPWR VPWR _16867_/Y sky130_fd_sc_hd__inv_2
X_19655_ _13251_/B VGND VGND VPWR VPWR _19655_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18377__D _14342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15818_ _15818_/A VGND VGND VPWR VPWR _15818_/X sky130_fd_sc_hd__buf_2
X_18606_ _24162_/Q VGND VGND VPWR VPWR _18606_/X sky130_fd_sc_hd__buf_2
X_19586_ _19586_/A VGND VGND VPWR VPWR _21694_/B sky130_fd_sc_hd__inv_2
X_16798_ _15019_/Y _16792_/X _16451_/X _16792_/X VGND VGND VPWR VPWR _16798_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_241_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22325__B2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18537_ _18537_/A VGND VGND VPWR VPWR _24183_/D sky130_fd_sc_hd__inv_2
XFILLER_206_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15749_ _15725_/A VGND VGND VPWR VPWR _15749_/X sky130_fd_sc_hd__buf_2
XFILLER_61_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18468_ _24179_/Q VGND VGND VPWR VPWR _18543_/A sky130_fd_sc_hd__inv_2
X_17419_ _17396_/A _17410_/A _24002_/Q _21008_/B _17413_/A VGND VGND VPWR VPWR _17419_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_221_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18399_ _16189_/Y _18490_/A _16189_/Y _18490_/A VGND VGND VPWR VPWR _18399_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12577__B1 _12618_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20430_ _20430_/A VGND VGND VPWR VPWR _20430_/X sky130_fd_sc_hd__buf_2
XFILLER_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17505__A1_N _25531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20361_ _20360_/Y _20352_/A _15656_/X _20352_/A VGND VGND VPWR VPWR _23420_/D sky130_fd_sc_hd__a2bb2o_4
X_22100_ _21277_/A _22076_/Y _22084_/Y _22092_/Y _22099_/Y VGND VGND VPWR VPWR _22100_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23080_ _24608_/Q _23189_/B VGND VGND VPWR VPWR _23080_/X sky130_fd_sc_hd__or2_4
XFILLER_161_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20292_ _21644_/B _20291_/X _16887_/X _20291_/X VGND VGND VPWR VPWR _20292_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22940__A _22940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_45_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22031_ _22034_/A _20369_/Y VGND VGND VPWR VPWR _22033_/B sky130_fd_sc_hd__or2_4
XFILLER_161_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21556__A _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17753__B _17753_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23945__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15554__A _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23982_ _24003_/CLK _21015_/Y HRESETn VGND VGND VPWR VPWR _21016_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_228_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22933_ _16003_/A VGND VGND VPWR VPWR _23140_/B sky130_fd_sc_hd__buf_2
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23108__A3 _22861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22864_ _22854_/B VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__buf_2
XANTENNA__22387__A _22387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24603_ _24989_/CLK _16418_/X HRESETn VGND VGND VPWR VPWR _24603_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21815_ _21815_/A _21815_/B _21815_/C VGND VGND VPWR VPWR _21815_/X sky130_fd_sc_hd__and3_4
X_22795_ _22787_/X _22791_/Y _22501_/X _22794_/X VGND VGND VPWR VPWR _22795_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16385__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24534_ _24566_/CLK _24534_/D HRESETn VGND VGND VPWR VPWR _24534_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21746_ _21565_/Y _21739_/X _21741_/X _21745_/Y VGND VGND VPWR VPWR _21746_/X sky130_fd_sc_hd__a211o_4
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _24430_/CLK _16774_/X HRESETn VGND VGND VPWR VPWR _22713_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21677_ _21485_/A _21677_/B _21677_/C VGND VGND VPWR VPWR _21677_/X sky130_fd_sc_hd__and3_4
XFILLER_196_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22834__B _23027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23684_/CLK _23416_/D VGND VGND VPWR VPWR _20372_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_11_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20628_ _17411_/X VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__buf_2
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24396_ _24407_/CLK _24396_/D HRESETn VGND VGND VPWR VPWR _16996_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15506__B1 HADDR[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20559_ _20559_/A VGND VGND VPWR VPWR _20559_/Y sky130_fd_sc_hd__inv_2
X_23347_ _16803_/A _22153_/X _22815_/X _23346_/X VGND VGND VPWR VPWR _23347_/X sky130_fd_sc_hd__a211o_4
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _13104_/A _13096_/X _13100_/C VGND VGND VPWR VPWR _25350_/D sky130_fd_sc_hd__and3_4
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14080_ _14063_/Y _14079_/X _14059_/X _14024_/X VGND VGND VPWR VPWR _14543_/B sky130_fd_sc_hd__or4_4
X_23278_ _22837_/X _23269_/Y _23273_/Y _23277_/X VGND VGND VPWR VPWR _23286_/C sky130_fd_sc_hd__a211o_4
XANTENNA__23044__A2 _22531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22850__A _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _12306_/A _13031_/B VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__or2_4
X_25017_ _25018_/CLK _25017_/D HRESETn VGND VGND VPWR VPWR _25017_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22229_ _22214_/A _22229_/B _22228_/X VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__or3_4
XFILLER_154_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21466__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_2_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17770_ _17761_/X _17770_/B VGND VGND VPWR VPWR _17770_/X sky130_fd_sc_hd__or2_4
X_14982_ _25035_/Q _14980_/Y _15075_/D _14978_/A VGND VGND VPWR VPWR _14982_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14493__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16721_ _16709_/A VGND VGND VPWR VPWR _16721_/X sky130_fd_sc_hd__buf_2
X_13933_ _24978_/Q VGND VGND VPWR VPWR _13933_/X sky130_fd_sc_hd__buf_2
XFILLER_208_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19440_ _19435_/Y _19438_/X _19439_/X _19438_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17431__B1 _17430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16652_ _16652_/A VGND VGND VPWR VPWR _16653_/A sky130_fd_sc_hd__inv_2
XFILLER_207_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13864_ _13872_/A VGND VGND VPWR VPWR _13864_/X sky130_fd_sc_hd__buf_2
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15603_ _15601_/Y _15597_/X _11797_/X _15602_/X VGND VGND VPWR VPWR _15603_/X sky130_fd_sc_hd__a2bb2o_4
X_12815_ _12815_/A VGND VGND VPWR VPWR _22678_/A sky130_fd_sc_hd__buf_2
X_19371_ _23771_/Q VGND VGND VPWR VPWR _19371_/Y sky130_fd_sc_hd__inv_2
X_16583_ _24539_/Q VGND VGND VPWR VPWR _16583_/Y sky130_fd_sc_hd__inv_2
X_13795_ _13795_/A VGND VGND VPWR VPWR _13795_/Y sky130_fd_sc_hd__inv_2
X_18322_ _18301_/X _18321_/Y _18302_/Y _18320_/X VGND VGND VPWR VPWR _18322_/X sky130_fd_sc_hd__o22a_4
X_15534_ _15532_/Y _15533_/X HADDR[9] _15533_/X VGND VGND VPWR VPWR _24939_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_203_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12746_ _12738_/B _12745_/X _12741_/C VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__and3_4
XFILLER_15_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18253_ _22595_/A _18243_/X _15761_/X _18252_/X VGND VGND VPWR VPWR _24242_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_203_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15465_ _15465_/A VGND VGND VPWR VPWR _20620_/A sky130_fd_sc_hd__buf_2
XANTENNA__15745__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12677_ _12676_/X VGND VGND VPWR VPWR _12678_/B sky130_fd_sc_hd__inv_2
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _16296_/A _24375_/Q _16296_/Y _17203_/Y VGND VGND VPWR VPWR _17204_/X sky130_fd_sc_hd__o22a_4
XFILLER_187_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _14415_/X VGND VGND VPWR VPWR _14416_/X sky130_fd_sc_hd__buf_2
XFILLER_147_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18184_ _17984_/A _18184_/B VGND VGND VPWR VPWR _18184_/X sky130_fd_sc_hd__or2_4
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15396_ _15396_/A _15299_/Y VGND VGND VPWR VPWR _15423_/B sky130_fd_sc_hd__or2_4
XFILLER_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15760__A3 _15759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17135_/A VGND VGND VPWR VPWR _17135_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14347_ _14347_/A VGND VGND VPWR VPWR _14347_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18865__A1_N _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17066_ _17060_/A _17059_/X _17062_/B _17065_/X VGND VGND VPWR VPWR _17067_/A sky130_fd_sc_hd__a211o_4
X_14278_ _14277_/Y _14273_/X _13809_/X _14273_/X VGND VGND VPWR VPWR _25193_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16170__B1 _15483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12274__A2_N _21715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16017_ _16016_/Y _16012_/X _15952_/X _16012_/X VGND VGND VPWR VPWR _24748_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13159__A _13212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13229_ _13385_/A _13229_/B VGND VGND VPWR VPWR _13229_/X sky130_fd_sc_hd__or2_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12063__A _21583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17968_ _17964_/X _17967_/X _18016_/A VGND VGND VPWR VPWR _17968_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _19706_/Y _19704_/X _19560_/X _19704_/X VGND VGND VPWR VPWR _19707_/X sky130_fd_sc_hd__a2bb2o_4
X_16919_ _24710_/Q _24287_/Q _16115_/Y _17753_/B VGND VGND VPWR VPWR _16922_/C sky130_fd_sc_hd__o22a_4
XANTENNA__13606__B _14442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17899_ _17899_/A VGND VGND VPWR VPWR _17913_/B sky130_fd_sc_hd__buf_2
XFILLER_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19638_ _19638_/A VGND VGND VPWR VPWR _19638_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14236__B1 _13846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19569_ _19568_/Y _19565_/X _19454_/X _19565_/X VGND VGND VPWR VPWR _23702_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15984__B1 _15905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21600_ _16723_/Y _22575_/A VGND VGND VPWR VPWR _21600_/X sky130_fd_sc_hd__and2_4
XFILLER_179_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22580_ _22768_/A _22580_/B VGND VGND VPWR VPWR _22580_/Y sky130_fd_sc_hd__nor2_4
XFILLER_178_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24694__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21531_ _21531_/A _23016_/A VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__or2_4
XANTENNA__15736__B1 _11776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23259__C1 _23258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24623__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21462_ _21461_/X VGND VGND VPWR VPWR _21528_/C sky130_fd_sc_hd__inv_2
X_24250_ _24252_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19478__B2 _19460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20413_ _20413_/A VGND VGND VPWR VPWR _20413_/Y sky130_fd_sc_hd__inv_2
X_23201_ _23118_/X _23201_/B VGND VGND VPWR VPWR _23208_/C sky130_fd_sc_hd__and2_4
XFILLER_147_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21393_ _14688_/X _19809_/Y VGND VGND VPWR VPWR _21393_/X sky130_fd_sc_hd__or2_4
X_24181_ _24523_/CLK _18546_/X HRESETn VGND VGND VPWR VPWR _24181_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12970__B1 _12875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20344_ _20343_/X VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__buf_2
X_23132_ _23208_/A _23132_/B _23132_/C _23131_/X VGND VGND VPWR VPWR _23132_/X sky130_fd_sc_hd__or4_4
XFILLER_146_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23063_ _22993_/X _23061_/X _23062_/X _25548_/Q _22793_/X VGND VGND VPWR VPWR _23063_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_161_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20275_ _20274_/Y _20270_/X _15656_/X _20270_/A VGND VGND VPWR VPWR _20275_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22014_ _13802_/A _21280_/A VGND VGND VPWR VPWR _22014_/X sky130_fd_sc_hd__or2_4
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18989__B1 _18969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_132_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23703_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23329__A3 _22145_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12701__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_195_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24657_/CLK sky130_fd_sc_hd__clkbuf_1
X_23965_ _23946_/CLK sda_i_S4 HRESETn VGND VGND VPWR VPWR _23966_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22916_ _21543_/A VGND VGND VPWR VPWR _23165_/B sky130_fd_sc_hd__buf_2
XFILLER_72_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23896_ _23880_/CLK _23896_/D VGND VGND VPWR VPWR _23896_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22847_ _23144_/A _22843_/X _22844_/X _22846_/X VGND VGND VPWR VPWR _22848_/A sky130_fd_sc_hd__o22a_4
XFILLER_25_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ _12599_/Y _24863_/Q _25407_/Q _12571_/Y VGND VGND VPWR VPWR _12607_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _13578_/A _14586_/C _13578_/Y _14590_/A VGND VGND VPWR VPWR _13580_/X sky130_fd_sc_hd__o22a_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22778_ _22778_/A _23322_/B VGND VGND VPWR VPWR _22778_/X sky130_fd_sc_hd__or2_4
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12531_ _12618_/B _24876_/Q _12529_/Y _24876_/Q VGND VGND VPWR VPWR _12531_/X sky130_fd_sc_hd__a2bb2o_4
X_24517_ _24684_/CLK _24517_/D HRESETn VGND VGND VPWR VPWR _24517_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21729_ _20610_/A _14203_/X _14472_/Y _17424_/X VGND VGND VPWR VPWR _21729_/X sky130_fd_sc_hd__o22a_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17939__A _18023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25497_ _24171_/CLK _12046_/X HRESETn VGND VGND VPWR VPWR _25497_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22564__B _21104_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15250_ _15250_/A _15249_/Y VGND VGND VPWR VPWR _15252_/B sky130_fd_sc_hd__or2_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12462_ _12464_/B VGND VGND VPWR VPWR _12462_/Y sky130_fd_sc_hd__inv_2
X_24448_ _25043_/CLK _16812_/X HRESETn VGND VGND VPWR VPWR _14939_/A sky130_fd_sc_hd__dfrtp_4
X_14201_ _14201_/A VGND VGND VPWR VPWR _21861_/A sky130_fd_sc_hd__buf_2
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15181_ _15081_/X _15181_/B VGND VGND VPWR VPWR _15181_/X sky130_fd_sc_hd__or2_4
X_12393_ _12393_/A _13017_/B VGND VGND VPWR VPWR _12394_/D sky130_fd_sc_hd__or2_4
X_24379_ _24378_/CLK _17172_/X HRESETn VGND VGND VPWR VPWR _17002_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14132_ _14131_/X _14132_/B VGND VGND VPWR VPWR _14133_/A sky130_fd_sc_hd__and2_4
X_14063_ _14063_/A VGND VGND VPWR VPWR _14063_/Y sky130_fd_sc_hd__inv_2
X_18940_ _18952_/A VGND VGND VPWR VPWR _18940_/X sky130_fd_sc_hd__buf_2
XFILLER_180_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13014_ _13014_/A _13011_/X VGND VGND VPWR VPWR _13014_/X sky130_fd_sc_hd__or2_4
XANTENNA__17393__B _17393_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18871_ _18867_/X _18868_/X _18869_/X _18871_/D VGND VGND VPWR VPWR _18872_/D sky130_fd_sc_hd__or4_4
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17822_ _17824_/B VGND VGND VPWR VPWR _17823_/B sky130_fd_sc_hd__inv_2
XANTENNA__16455__B2 _16384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14466__B1 _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12611__A _12638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21924__A _22093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14965_ _14965_/A VGND VGND VPWR VPWR _15079_/A sky130_fd_sc_hd__buf_2
X_17753_ _17753_/A _17753_/B VGND VGND VPWR VPWR _17753_/X sky130_fd_sc_hd__or2_4
XFILLER_207_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13916_ _13916_/A VGND VGND VPWR VPWR _13916_/Y sky130_fd_sc_hd__inv_2
X_16704_ _16709_/A VGND VGND VPWR VPWR _16704_/X sky130_fd_sc_hd__buf_2
X_17684_ _17684_/A _17684_/B VGND VGND VPWR VPWR _17685_/C sky130_fd_sc_hd__nand2_4
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14896_ _14895_/X _16845_/A _14895_/X _16845_/A VGND VGND VPWR VPWR _14905_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21751__A2 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16635_ RsRx_S0 _16182_/B _16634_/Y VGND VGND VPWR VPWR _16643_/B sky130_fd_sc_hd__o21a_4
X_19423_ _19420_/Y _19415_/X _19421_/X _19422_/X VGND VGND VPWR VPWR _19423_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13847_ _13560_/Y _13842_/X _13846_/X _13842_/X VGND VGND VPWR VPWR _13847_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15966__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19157__B1 _19131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16566_ _16566_/A VGND VGND VPWR VPWR _16566_/Y sky130_fd_sc_hd__inv_2
X_19354_ _19352_/Y _19348_/X _19308_/X _19353_/X VGND VGND VPWR VPWR _19354_/X sky130_fd_sc_hd__a2bb2o_4
X_13778_ _13778_/A VGND VGND VPWR VPWR _14611_/A sky130_fd_sc_hd__inv_2
XFILLER_200_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22755__A _22755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15981__A3 _16248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15517_ _15517_/A VGND VGND VPWR VPWR _15517_/Y sky130_fd_sc_hd__inv_2
X_18305_ _18301_/A VGND VGND VPWR VPWR _18306_/A sky130_fd_sc_hd__buf_2
XANTENNA__22700__B2 _22289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12729_ _12729_/A _12713_/X VGND VGND VPWR VPWR _12729_/Y sky130_fd_sc_hd__nand2_4
X_19285_ _19285_/A VGND VGND VPWR VPWR _22077_/B sky130_fd_sc_hd__inv_2
X_16497_ _24572_/Q VGND VGND VPWR VPWR _16497_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18236_ _15703_/X _18220_/X _18235_/X _24248_/Q _18029_/A VGND VGND VPWR VPWR _18236_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_148_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15448_ _13933_/X _15446_/X _15441_/X _24979_/Q _15447_/X VGND VGND VPWR VPWR _15448_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23256__A2 _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15733__A3 _15732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _18199_/A _23831_/Q VGND VGND VPWR VPWR _18169_/B sky130_fd_sc_hd__or2_4
XFILLER_191_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15379_ _15384_/A _15376_/B _15378_/Y VGND VGND VPWR VPWR _24998_/D sky130_fd_sc_hd__and3_4
XFILLER_156_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17118_ _17118_/A _17115_/B VGND VGND VPWR VPWR _17119_/C sky130_fd_sc_hd__nand2_4
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18098_ _18098_/A VGND VGND VPWR VPWR _18164_/A sky130_fd_sc_hd__buf_2
X_17049_ _24389_/Q VGND VGND VPWR VPWR _17050_/C sky130_fd_sc_hd__inv_2
XFILLER_131_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20060_ _20059_/Y VGND VGND VPWR VPWR _20060_/X sky130_fd_sc_hd__buf_2
XANTENNA__15815__A1_N _12330_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_205_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24556_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21990__A2 _20360_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21834__A _21834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23192__A1 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22649__B _23053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23750_ _23735_/CLK _23750_/D VGND VGND VPWR VPWR _18181_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16452__A2_N _16446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20962_ _20960_/Y _20957_/X _20961_/X VGND VGND VPWR VPWR _20962_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22701_ _23144_/A VGND VGND VPWR VPWR _23008_/A sky130_fd_sc_hd__buf_2
XANTENNA__24875__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23799_/CLK _19637_/X VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _20891_/Y _20888_/Y _20896_/A VGND VGND VPWR VPWR _20893_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25420_ _25425_/CLK _12700_/Y HRESETn VGND VGND VPWR VPWR _25420_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24804__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22632_ _22523_/X _22630_/X _21968_/X _22631_/Y VGND VGND VPWR VPWR _22632_/X sky130_fd_sc_hd__o22a_4
XFILLER_159_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25351_ _25368_/CLK _13098_/X HRESETn VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__dfrtp_4
X_22563_ _22562_/X VGND VGND VPWR VPWR _22563_/X sky130_fd_sc_hd__buf_2
XANTENNA__20702__B1 _20698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24302_ _24302_/CLK _17692_/X HRESETn VGND VGND VPWR VPWR _17504_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21514_ _21514_/A _21282_/X VGND VGND VPWR VPWR _21514_/X sky130_fd_sc_hd__or2_4
X_25282_ _23516_/CLK _13777_/X HRESETn VGND VGND VPWR VPWR _25282_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22494_ _22721_/B VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__buf_2
XFILLER_166_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15724__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24233_ _24233_/CLK _24233_/D HRESETn VGND VGND VPWR VPWR _24233_/Q sky130_fd_sc_hd__dfrtp_4
X_21445_ _22202_/C VGND VGND VPWR VPWR _21445_/X sky130_fd_sc_hd__buf_2
XFILLER_194_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21376_ _14221_/Y _14202_/X _14282_/Y _21375_/X VGND VGND VPWR VPWR _21377_/D sky130_fd_sc_hd__o22a_4
X_24164_ _25145_/CLK _18601_/X HRESETn VGND VGND VPWR VPWR _24164_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20327_ _22253_/B _20324_/X _19993_/X _20324_/X VGND VGND VPWR VPWR _23434_/D sky130_fd_sc_hd__a2bb2o_4
X_23115_ _21316_/X VGND VGND VPWR VPWR _23115_/X sky130_fd_sc_hd__buf_2
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24095_ _24095_/CLK _20546_/X HRESETn VGND VGND VPWR VPWR _24095_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20258_ _20270_/A VGND VGND VPWR VPWR _20258_/X sky130_fd_sc_hd__buf_2
X_23046_ _23045_/X VGND VGND VPWR VPWR _23046_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20189_ _20188_/Y _20184_/X _20146_/X _20172_/A VGND VGND VPWR VPWR _20189_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24997_ _24981_/CLK _24997_/D HRESETn VGND VGND VPWR VPWR _15092_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14750_ _14731_/X _14738_/Y _14749_/X _22055_/A _14732_/Y VGND VGND VPWR VPWR _25071_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11962_ _11960_/Y _11956_/X _11961_/X _11956_/X VGND VGND VPWR VPWR _25509_/D sky130_fd_sc_hd__a2bb2o_4
X_23948_ _23395_/CLK _20994_/A HRESETn VGND VGND VPWR VPWR _20996_/C sky130_fd_sc_hd__dfstp_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_1_HCLK clkbuf_1_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_245_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13701_ _13707_/B VGND VGND VPWR VPWR _13702_/B sky130_fd_sc_hd__inv_2
X_14681_ _19166_/A _19166_/B _19166_/A _19166_/B VGND VGND VPWR VPWR _25077_/D sky130_fd_sc_hd__a2bb2o_4
X_11893_ _11892_/Y _11887_/B VGND VGND VPWR VPWR _11893_/X sky130_fd_sc_hd__and2_4
X_23879_ _23459_/CLK _19069_/X VGND VGND VPWR VPWR _19067_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_205_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16420_ _15131_/Y _16415_/X _16419_/X _16415_/X VGND VGND VPWR VPWR _24602_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _14801_/B VGND VGND VPWR VPWR _13636_/C sky130_fd_sc_hd__inv_2
XFILLER_71_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22575__A _22575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16351_ _24626_/Q VGND VGND VPWR VPWR _16351_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13563_ _13563_/A _13556_/X _13563_/C _13563_/D VGND VGND VPWR VPWR _13597_/A sky130_fd_sc_hd__or4_4
X_25549_ _25539_/CLK _25549_/D HRESETn VGND VGND VPWR VPWR _25549_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15302_ _25009_/Q VGND VGND VPWR VPWR _15302_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12514_ _12514_/A _12514_/B _12513_/Y VGND VGND VPWR VPWR _25439_/D sky130_fd_sc_hd__and3_4
X_19070_ _23878_/Q VGND VGND VPWR VPWR _19070_/Y sky130_fd_sc_hd__inv_2
X_16282_ _15667_/A _16001_/X VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__or2_4
X_13494_ _13493_/Y _13491_/X _11856_/X _13491_/X VGND VGND VPWR VPWR _13494_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16373__B1 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18021_ _18129_/A _23843_/Q VGND VGND VPWR VPWR _18021_/X sky130_fd_sc_hd__or2_4
X_15233_ _14921_/X _15232_/X VGND VGND VPWR VPWR _15234_/C sky130_fd_sc_hd__nand2_4
X_12445_ _12293_/Y _12442_/X VGND VGND VPWR VPWR _12445_/X sky130_fd_sc_hd__or2_4
XFILLER_173_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15164_ _25011_/Q VGND VGND VPWR VPWR _15164_/Y sky130_fd_sc_hd__inv_2
X_12376_ _13026_/A _24851_/Q _25360_/Q _12375_/Y VGND VGND VPWR VPWR _12380_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22461__A3 _16468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14115_ _14128_/C _14115_/B _14114_/Y VGND VGND VPWR VPWR _14115_/X sky130_fd_sc_hd__and3_4
XFILLER_126_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15095_ _15095_/A VGND VGND VPWR VPWR _15095_/Y sky130_fd_sc_hd__inv_2
X_19972_ _19979_/A VGND VGND VPWR VPWR _19972_/X sky130_fd_sc_hd__buf_2
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22749__A1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14046_ _14062_/A _14008_/X _14062_/C VGND VGND VPWR VPWR _14047_/A sky130_fd_sc_hd__or3_4
X_18923_ _22080_/B _18917_/X _16881_/X _18922_/X VGND VGND VPWR VPWR _23930_/D sky130_fd_sc_hd__a2bb2o_4
X_18854_ _24556_/Q _18685_/Y _16532_/A _18810_/A VGND VGND VPWR VPWR _18854_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17805_ _17807_/B VGND VGND VPWR VPWR _17805_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15997_ _12240_/Y _15990_/X _15848_/X _15947_/A VGND VGND VPWR VPWR _15997_/X sky130_fd_sc_hd__a2bb2o_4
X_18785_ _18699_/B _18779_/X _18740_/X _18782_/B VGND VGND VPWR VPWR _18786_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16748__A _16762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19378__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23174__B2 _22924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14948_ _14937_/X _14940_/X _14948_/C _14947_/X VGND VGND VPWR VPWR _14948_/X sky130_fd_sc_hd__or4_4
X_17736_ _17732_/X _17735_/X _17732_/X _17735_/X VGND VGND VPWR VPWR _17736_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_35_0_HCLK clkbuf_8_34_0_HCLK/A VGND VGND VPWR VPWR _25068_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20070__A2_N _20065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14879_ _14889_/A _24006_/Q VGND VGND VPWR VPWR _14879_/X sky130_fd_sc_hd__or2_4
X_17667_ _17667_/A _17667_/B VGND VGND VPWR VPWR _17668_/C sky130_fd_sc_hd__or2_4
Xclkbuf_8_98_0_HCLK clkbuf_7_49_0_HCLK/X VGND VGND VPWR VPWR _24641_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _19404_/Y _19405_/X _19383_/X _19405_/X VGND VGND VPWR VPWR _23759_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16618_ _16618_/A VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__buf_2
XFILLER_23_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17598_ _17598_/A _17598_/B _17597_/Y VGND VGND VPWR VPWR _24327_/D sky130_fd_sc_hd__and3_4
XFILLER_210_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _16548_/Y _16469_/X _16375_/X _16469_/X VGND VGND VPWR VPWR _24552_/D sky130_fd_sc_hd__a2bb2o_4
X_19337_ _23783_/Q VGND VGND VPWR VPWR _19337_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22685__B1 _21591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16483__A _16495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19268_ _23808_/Q VGND VGND VPWR VPWR _19268_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ _18059_/A _18215_/X _18218_/X VGND VGND VPWR VPWR _18220_/C sky130_fd_sc_hd__or3_4
X_19199_ _19198_/Y _19196_/X _19085_/X _19196_/X VGND VGND VPWR VPWR _23833_/D sky130_fd_sc_hd__a2bb2o_4
X_21230_ _21032_/X VGND VGND VPWR VPWR _21868_/B sky130_fd_sc_hd__buf_2
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21161_ _21161_/A VGND VGND VPWR VPWR _21161_/X sky130_fd_sc_hd__buf_2
XFILLER_160_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17745__C _21834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20112_ _24415_/Q VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__buf_2
XFILLER_236_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21092_ _21023_/B _21105_/B VGND VGND VPWR VPWR _21092_/X sky130_fd_sc_hd__and2_4
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20043_ _20043_/A VGND VGND VPWR VPWR _20043_/Y sky130_fd_sc_hd__inv_2
X_24920_ _24029_/CLK _15593_/X HRESETn VGND VGND VPWR VPWR _15592_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_219_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24851_ _24889_/CLK _15813_/X HRESETn VGND VGND VPWR VPWR _24851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22328__A1_N _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23802_ _23514_/CLK _19287_/X VGND VGND VPWR VPWR _19285_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15562__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24782_ _24792_/CLK _24782_/D HRESETn VGND VGND VPWR VPWR _24782_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21176__B1 _16379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _18366_/Y _21995_/B _18355_/Y _23422_/Q VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__o22a_4
XPHY_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23733_ _23735_/CLK _23733_/D VGND VGND VPWR VPWR _19477_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_121_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _20943_/Y _20940_/Y _20949_/B VGND VGND VPWR VPWR _20945_/X sky130_fd_sc_hd__o21a_4
XPHY_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23654_/CLK _23664_/D VGND VGND VPWR VPWR _13361_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_198_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_6_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _16706_/Y _20854_/X _20863_/X _20875_/X VGND VGND VPWR VPWR _20876_/X sky130_fd_sc_hd__o22a_4
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25403_ _24799_/CLK _25403_/D HRESETn VGND VGND VPWR VPWR _25403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22615_ _15618_/Y _22577_/B VGND VGND VPWR VPWR _22615_/X sky130_fd_sc_hd__and2_4
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _23563_/CLK _23595_/D VGND VGND VPWR VPWR _23595_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16393__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25334_ _25488_/CLK _13377_/X HRESETn VGND VGND VPWR VPWR _25334_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22546_ _15032_/A _22543_/X _22545_/X VGND VGND VPWR VPWR _22546_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16355__B1 _16157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25265_ _25309_/CLK _13850_/X HRESETn VGND VGND VPWR VPWR _25265_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22477_ _22298_/X VGND VGND VPWR VPWR _22479_/A sky130_fd_sc_hd__buf_2
X_12230_ _22483_/A VGND VGND VPWR VPWR _12230_/Y sky130_fd_sc_hd__inv_2
X_24216_ _25292_/CLK _18328_/X HRESETn VGND VGND VPWR VPWR _21834_/A sky130_fd_sc_hd__dfstp_4
XFILLER_5_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21428_ _21029_/A VGND VGND VPWR VPWR _21535_/A sky130_fd_sc_hd__buf_2
XANTENNA__16107__B1 _15950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25196_ _25200_/CLK _14271_/X HRESETn VGND VGND VPWR VPWR _14270_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21100__B1 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12161_ _24120_/Q VGND VGND VPWR VPWR _12161_/Y sky130_fd_sc_hd__inv_2
X_24147_ _24145_/CLK _24147_/D HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_21359_ _14406_/Y _14202_/X _14499_/Y _14266_/A VGND VGND VPWR VPWR _21359_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12092_ _12092_/A VGND VGND VPWR VPWR _12092_/Y sky130_fd_sc_hd__inv_2
X_24078_ _24029_/CLK _24078_/D HRESETn VGND VGND VPWR VPWR _13677_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13257__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15920_ _13548_/A _15920_/B VGND VGND VPWR VPWR _15922_/A sky130_fd_sc_hd__or2_4
X_23029_ _22836_/A _23029_/B _23029_/C VGND VGND VPWR VPWR _23029_/X sky130_fd_sc_hd__and3_4
XANTENNA__18649__A1_N _24521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25140__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13892__A1 _24007_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15851_ _19761_/A VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__buf_2
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24797__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14802_ _14801_/X VGND VGND VPWR VPWR _14802_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24726__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15782_ _19761_/A VGND VGND VPWR VPWR _15782_/X sky130_fd_sc_hd__buf_2
X_18570_ _18418_/Y _18569_/X VGND VGND VPWR VPWR _18570_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_251_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _24343_/CLK sky130_fd_sc_hd__clkbuf_1
X_12994_ _12994_/A VGND VGND VPWR VPWR _13021_/A sky130_fd_sc_hd__inv_2
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14901__A1_N _25019_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14733_ _14712_/A _14713_/A _14729_/Y _13748_/A _14732_/Y VGND VGND VPWR VPWR _14733_/X
+ sky130_fd_sc_hd__a32o_4
X_17521_ _25549_/Q _24320_/Q _11775_/Y _17520_/Y VGND VGND VPWR VPWR _17521_/X sky130_fd_sc_hd__o22a_4
X_11945_ _11942_/Y _11935_/X _11943_/X _11944_/X VGND VGND VPWR VPWR _11945_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _19139_/A VGND VGND VPWR VPWR _17452_/X sky130_fd_sc_hd__buf_2
XANTENNA__16912__A2_N _21066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14664_ _17950_/A _14650_/C _14662_/X VGND VGND VPWR VPWR _25080_/D sky130_fd_sc_hd__o21a_4
XFILLER_221_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11876_ _13481_/A VGND VGND VPWR VPWR _11876_/X sky130_fd_sc_hd__buf_2
X_16403_ _16415_/A VGND VGND VPWR VPWR _16403_/X sky130_fd_sc_hd__buf_2
X_13615_ _13615_/A VGND VGND VPWR VPWR _13615_/Y sky130_fd_sc_hd__inv_2
X_17383_ _17357_/A _17356_/X _17298_/A _17380_/Y VGND VGND VPWR VPWR _17384_/A sky130_fd_sc_hd__a211o_4
XFILLER_189_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14595_ _14595_/A VGND VGND VPWR VPWR _14595_/X sky130_fd_sc_hd__buf_2
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14816__A _14816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16334_ HWDATA[16] VGND VGND VPWR VPWR _16334_/X sky130_fd_sc_hd__buf_2
X_19122_ _19118_/Y _19121_/X _19032_/X _19121_/X VGND VGND VPWR VPWR _23860_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16734__C _22592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13546_ _13652_/A _13543_/Y _13481_/X _13543_/Y VGND VGND VPWR VPWR _25308_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_197_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15149__B2 _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20142__B2 _20141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19053_ _13634_/X VGND VGND VPWR VPWR _19143_/B sky130_fd_sc_hd__buf_2
XFILLER_185_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16265_ _16263_/Y _16264_/X _16070_/X _16264_/X VGND VGND VPWR VPWR _24658_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22419__B1 _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13477_ _21577_/B VGND VGND VPWR VPWR _13504_/B sky130_fd_sc_hd__buf_2
XFILLER_127_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _15215_/X VGND VGND VPWR VPWR _25035_/D sky130_fd_sc_hd__inv_2
X_18004_ _17954_/A _17989_/X _18004_/C VGND VGND VPWR VPWR _18004_/X sky130_fd_sc_hd__and3_4
XFILLER_127_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12428_ _12428_/A _12428_/B VGND VGND VPWR VPWR _12429_/C sky130_fd_sc_hd__or2_4
XANTENNA__19854__A2_N _19851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16196_ _16202_/A VGND VGND VPWR VPWR _16196_/X sky130_fd_sc_hd__buf_2
X_15147_ _15306_/B _24602_/Q _25002_/Q _15098_/Y VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24342__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ _12997_/D _24839_/Q _12997_/D _24839_/Q VGND VGND VPWR VPWR _12360_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21368__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18023__A _18023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23286__D _23285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12183__A1_N SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15078_ _15073_/X _15078_/B VGND VGND VPWR VPWR _15078_/X sky130_fd_sc_hd__or2_4
X_19955_ _23568_/Q VGND VGND VPWR VPWR _19955_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14029_ _14545_/A _14028_/X VGND VGND VPWR VPWR _14029_/Y sky130_fd_sc_hd__nand2_4
X_18906_ _18905_/X VGND VGND VPWR VPWR _20430_/A sky130_fd_sc_hd__inv_2
X_19886_ _19885_/Y _19883_/X _19629_/X _19883_/X VGND VGND VPWR VPWR _23595_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_61_0_HCLK clkbuf_5_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18271__B1 _16791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18837_ _16548_/Y _18621_/X _16548_/Y _18621_/X VGND VGND VPWR VPWR _18837_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22199__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18768_ _18768_/A _18768_/B VGND VGND VPWR VPWR _18769_/C sky130_fd_sc_hd__or2_4
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17719_ _24221_/Q VGND VGND VPWR VPWR _18289_/C sky130_fd_sc_hd__inv_2
XANTENNA__19789__A _19788_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18699_ _18699_/A _18699_/B _18699_/C _18752_/A VGND VGND VPWR VPWR _18700_/B sky130_fd_sc_hd__or4_4
XFILLER_208_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20730_ _20730_/A VGND VGND VPWR VPWR _20730_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16585__B1 _16414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20661_ _20661_/A _20660_/Y _20669_/C VGND VGND VPWR VPWR _20661_/X sky130_fd_sc_hd__and3_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22122__A2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22400_ _22400_/A _22399_/Y VGND VGND VPWR VPWR _22401_/D sky130_fd_sc_hd__nor2_4
XANTENNA__12071__B1 _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20592_ _23958_/Q _18885_/B VGND VGND VPWR VPWR _20592_/Y sky130_fd_sc_hd__nand2_4
X_23380_ _21023_/X VGND VGND VPWR VPWR IRQ[24] sky130_fd_sc_hd__buf_2
XANTENNA__16337__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14445__B _14388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22331_ _12140_/A _12107_/A _18376_/Y _12080_/A VGND VGND VPWR VPWR _22331_/X sky130_fd_sc_hd__o22a_4
XFILLER_177_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22662__B _22662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25050_ _24000_/CLK _25050_/D HRESETn VGND VGND VPWR VPWR _14822_/C sky130_fd_sc_hd__dfrtp_4
X_22262_ _21685_/X _22262_/B _22261_/X VGND VGND VPWR VPWR _22262_/X sky130_fd_sc_hd__and3_4
XANTENNA__21559__A _21351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24001_ _24340_/CLK scl_i_S5 HRESETn VGND VGND VPWR VPWR _24002_/D sky130_fd_sc_hd__dfrtp_4
X_21213_ _21209_/X _21212_/X _24219_/Q VGND VGND VPWR VPWR _21213_/X sky130_fd_sc_hd__o21a_4
XFILLER_151_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22193_ _14270_/Y _14266_/A _17429_/Y _17424_/A VGND VGND VPWR VPWR _22193_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14461__A _14116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21144_ _21348_/B _21143_/X _17450_/B VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__o21a_4
XFILLER_160_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21075_ _21022_/B _21109_/B VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__and2_4
XFILLER_58_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24127__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20026_ _23544_/Q VGND VGND VPWR VPWR _21811_/B sky130_fd_sc_hd__inv_2
X_24903_ _24020_/CLK _24903_/D HRESETn VGND VGND VPWR VPWR _15634_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21294__A _21122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24890__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17491__B _17459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15292__A _15292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24834_ _24849_/CLK _15837_/X HRESETn VGND VGND VPWR VPWR _24834_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15001__A1_N _15292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24765_ _24765_/CLK _24765_/D HRESETn VGND VGND VPWR VPWR _22644_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19699__A _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21977_ _14635_/Y _19610_/A _25086_/Q _19614_/Y VGND VGND VPWR VPWR _21977_/X sky130_fd_sc_hd__o22a_4
XPHY_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19762__B1 _19761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11729_/X VGND VGND VPWR VPWR _11730_/Y sky130_fd_sc_hd__inv_2
X_23716_ _23716_/CLK _23716_/D VGND VGND VPWR VPWR _23716_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _13659_/A VGND VGND VPWR VPWR _20928_/Y sky130_fd_sc_hd__inv_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24696_ _24697_/CLK _16151_/X HRESETn VGND VGND VPWR VPWR _22574_/A sky130_fd_sc_hd__dfrtp_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_81_0_HCLK clkbuf_7_40_0_HCLK/X VGND VGND VPWR VPWR _25392_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15918__A3 _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/A _11979_/C VGND VGND VPWR VPWR _11661_/X sky130_fd_sc_hd__and2_4
X_23647_ _23647_/CLK _23647_/D VGND VGND VPWR VPWR _13400_/B sky130_fd_sc_hd__dfxtp_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20859_ _20865_/B VGND VGND VPWR VPWR _20859_/Y sky130_fd_sc_hd__inv_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18317__A1 _21676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13243_/X _13400_/B VGND VGND VPWR VPWR _13400_/X sky130_fd_sc_hd__or2_4
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _14364_/A _14379_/X _12097_/A _14369_/A VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16328__B1 _15970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23578_ _23514_/CLK _19932_/X VGND VGND VPWR VPWR _19930_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _13241_/X _13327_/X _13331_/C VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__or3_4
X_25317_ _25188_/CLK _25317_/D HRESETn VGND VGND VPWR VPWR _13514_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22529_ _22529_/A _22528_/X VGND VGND VPWR VPWR _22529_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_2_1_0_HCLK clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _16048_/Y _16044_/X _11813_/X _16049_/X VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13262_ _13372_/A _19819_/A VGND VGND VPWR VPWR _13263_/C sky130_fd_sc_hd__or2_4
X_25248_ _24003_/CLK _13982_/X HRESETn VGND VGND VPWR VPWR scl_oen_o_S5 sky130_fd_sc_hd__dfstp_4
X_15001_ _15292_/A _24452_/Q _15282_/A _15000_/Y VGND VGND VPWR VPWR _15005_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12213_ _12213_/A VGND VGND VPWR VPWR _12213_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13193_ _13197_/A _13193_/B _13193_/C VGND VGND VPWR VPWR _13193_/X sky130_fd_sc_hd__and3_4
X_25179_ _25181_/CLK _14327_/X HRESETn VGND VGND VPWR VPWR _25179_/Q sky130_fd_sc_hd__dfrtp_4
X_12144_ _12122_/A _12142_/X _12122_/Y _12143_/Y VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19740_ _13175_/B VGND VGND VPWR VPWR _19740_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24907__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12075_ _21577_/A VGND VGND VPWR VPWR _12109_/C sky130_fd_sc_hd__buf_2
X_16952_ _24285_/Q VGND VGND VPWR VPWR _16952_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15903_ _15714_/X _15902_/X _16252_/A _22605_/A _15871_/X VGND VGND VPWR VPWR _15903_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18253__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19671_ _13461_/B VGND VGND VPWR VPWR _19671_/Y sky130_fd_sc_hd__inv_2
X_16883_ _20115_/A VGND VGND VPWR VPWR _19803_/A sky130_fd_sc_hd__buf_2
XFILLER_77_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24560__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ _21167_/A _18621_/X _21167_/A _18621_/X VGND VGND VPWR VPWR _18622_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15834_ _15833_/X _15828_/X _16252_/A _24836_/Q _15802_/A VGND VGND VPWR VPWR _15834_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18553_ _18550_/A _18543_/B _18552_/X VGND VGND VPWR VPWR _18553_/X sky130_fd_sc_hd__and3_4
XANTENNA__22888__B1 _12773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12977_ _12828_/X _12950_/X _12891_/X _12974_/Y VGND VGND VPWR VPWR _12978_/A sky130_fd_sc_hd__a211o_4
X_15765_ HWDATA[9] VGND VGND VPWR VPWR _15765_/X sky130_fd_sc_hd__buf_2
XFILLER_80_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17504_ _17504_/A VGND VGND VPWR VPWR _17504_/Y sky130_fd_sc_hd__inv_2
X_11928_ _11910_/X _11919_/X VGND VGND VPWR VPWR _11928_/Y sky130_fd_sc_hd__nor2_4
X_14716_ _14715_/X VGND VGND VPWR VPWR _14716_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19402__A _19131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15696_ _15696_/A _15696_/B _15696_/C VGND VGND VPWR VPWR _15696_/X sky130_fd_sc_hd__or3_4
X_18484_ _18474_/Y _18484_/B _18557_/B VGND VGND VPWR VPWR _18515_/B sky130_fd_sc_hd__or3_4
X_14647_ _13547_/Y _13610_/X _13644_/A VGND VGND VPWR VPWR _14650_/C sky130_fd_sc_hd__o21a_4
X_17435_ _17432_/Y _17426_/X _17433_/X _17434_/X VGND VGND VPWR VPWR _17435_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11859_ _25528_/Q VGND VGND VPWR VPWR _11859_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_109_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24029_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18018__A _18098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__A2 _22299_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ _14577_/X VGND VGND VPWR VPWR _14578_/Y sky130_fd_sc_hd__inv_2
X_17366_ _17366_/A VGND VGND VPWR VPWR _24356_/D sky130_fd_sc_hd__inv_2
XFILLER_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19105_ _19099_/Y VGND VGND VPWR VPWR _19105_/X sky130_fd_sc_hd__buf_2
X_13529_ _13529_/A VGND VGND VPWR VPWR _20972_/B sky130_fd_sc_hd__buf_2
X_16317_ _16317_/A VGND VGND VPWR VPWR _16317_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17297_ _17267_/B _17276_/X _17245_/Y VGND VGND VPWR VPWR _17297_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16248_ _16248_/A VGND VGND VPWR VPWR _16248_/X sky130_fd_sc_hd__buf_2
X_19036_ _23890_/Q VGND VGND VPWR VPWR _19036_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19808__B2 _19806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16179_ _16179_/A VGND VGND VPWR VPWR _16179_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15845__A2 _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24648__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19938_ _19925_/Y VGND VGND VPWR VPWR _19938_/X sky130_fd_sc_hd__buf_2
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21379__B1 _21367_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18244__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _23601_/Q VGND VGND VPWR VPWR _21917_/B sky130_fd_sc_hd__inv_2
XFILLER_110_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22003__A _22003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21900_ _21895_/X _21900_/B VGND VGND VPWR VPWR _21900_/X sky130_fd_sc_hd__or2_4
XANTENNA__13625__A _18102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22880_ _22880_/A VGND VGND VPWR VPWR _22880_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16001__A _14199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22938__A _23008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21831_ _21827_/X _21830_/X _21697_/X VGND VGND VPWR VPWR _21831_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24550_ _24562_/CLK _24550_/D HRESETn VGND VGND VPWR VPWR _24550_/Q sky130_fd_sc_hd__dfrtp_4
X_21762_ _21731_/Y _21746_/X _21762_/C _21761_/X VGND VGND VPWR VPWR _21762_/X sky130_fd_sc_hd__or4_4
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_68_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_68_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23501_ _23690_/CLK _20147_/X VGND VGND VPWR VPWR _20145_/A sky130_fd_sc_hd__dfxtp_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20713_ _13135_/A _13134_/X _20712_/Y VGND VGND VPWR VPWR _20713_/Y sky130_fd_sc_hd__a21oi_4
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24481_ _25043_/CLK _16741_/X HRESETn VGND VGND VPWR VPWR _15026_/A sky130_fd_sc_hd__dfrtp_4
X_21693_ _21808_/A _21691_/X _21692_/X VGND VGND VPWR VPWR _21693_/X sky130_fd_sc_hd__and3_4
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23432_ _23553_/CLK _20332_/X VGND VGND VPWR VPWR _20331_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20644_ _15474_/Y _20623_/X _20637_/X _20643_/X VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__a211o_4
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23363_ _11979_/C _11970_/D _11968_/X VGND VGND VPWR VPWR _25558_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__17767__A _17767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20575_ _18881_/A _20571_/A VGND VGND VPWR VPWR _20575_/Y sky130_fd_sc_hd__nand2_4
XFILLER_137_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25102_ _25103_/CLK _25102_/D HRESETn VGND VGND VPWR VPWR _25102_/Q sky130_fd_sc_hd__dfrtp_4
X_22314_ _16615_/A _21330_/X _21331_/X _22313_/X VGND VGND VPWR VPWR _22315_/C sky130_fd_sc_hd__a211o_4
X_23294_ _23124_/X _23293_/X _21532_/X _16008_/A _21538_/X VGND VGND VPWR VPWR _23295_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16730__B1 _16729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17486__B _17459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25033_ _25030_/CLK _25033_/D HRESETn VGND VGND VPWR VPWR _25033_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13544__B1 _13524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22245_ _22027_/A _22245_/B VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__or2_4
XFILLER_127_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22176_ _14395_/Y _22176_/B VGND VGND VPWR VPWR _22183_/A sky130_fd_sc_hd__nor2_4
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21127_ _21025_/B _16280_/A _15663_/X _23386_/D _15667_/A VGND VGND VPWR VPWR _21127_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21058_ _21058_/A _21044_/X _21058_/C VGND VGND VPWR VPWR _21058_/X sky130_fd_sc_hd__and3_4
XANTENNA__11858__B1 _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _12850_/A _12900_/B VGND VGND VPWR VPWR _12901_/C sky130_fd_sc_hd__or2_4
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20009_ _20009_/A VGND VGND VPWR VPWR _21497_/B sky130_fd_sc_hd__inv_2
XFILLER_247_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13880_ _24007_/Q VGND VGND VPWR VPWR _13880_/X sky130_fd_sc_hd__buf_2
XANTENNA__16797__B1 _16796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ _24810_/Q VGND VGND VPWR VPWR _12831_/Y sky130_fd_sc_hd__inv_2
X_24817_ _24803_/CLK _15881_/X HRESETn VGND VGND VPWR VPWR _23199_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21843__A2_N _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19735__B1 _19734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15550_ _15549_/Y _15547_/X HADDR[1] _15547_/X VGND VGND VPWR VPWR _24931_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12762_ _12762_/A VGND VGND VPWR VPWR _12921_/C sky130_fd_sc_hd__buf_2
X_24748_ _24642_/CLK _24748_/D HRESETn VGND VGND VPWR VPWR _24748_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16549__B1 _16375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _25119_/Q VGND VGND VPWR VPWR _14501_/Y sky130_fd_sc_hd__inv_2
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A VGND VGND VPWR VPWR _11713_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15479_/Y _15477_/X _15480_/X _15477_/X VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_199_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12680_/A _12689_/X _12693_/C VGND VGND VPWR VPWR _12693_/X sky130_fd_sc_hd__and3_4
X_24679_ _24657_/CLK _16208_/X HRESETn VGND VGND VPWR VPWR _23218_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _25146_/Q VGND VGND VPWR VPWR _14432_/Y sky130_fd_sc_hd__inv_2
X_17220_ _17213_/X _17220_/B _17218_/X _17219_/X VGND VGND VPWR VPWR _17239_/A sky130_fd_sc_hd__or4_4
XFILLER_203_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22583__A _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _17142_/A _17142_/B VGND VGND VPWR VPWR _17152_/C sky130_fd_sc_hd__nand2_4
XANTENNA__12586__B2 _24875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _14369_/A VGND VGND VPWR VPWR _14364_/A sky130_fd_sc_hd__inv_2
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16581__A _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _24715_/Q VGND VGND VPWR VPWR _16102_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13310_/X _13312_/X _13313_/X VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__and3_4
X_17082_ _17095_/A _17082_/B _17081_/X VGND VGND VPWR VPWR _24405_/D sky130_fd_sc_hd__and3_4
X_14294_ _23444_/Q _14289_/X _14293_/A _25189_/Q _14293_/Y VGND VGND VPWR VPWR _25189_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16033_ _24741_/Q VGND VGND VPWR VPWR _16033_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12338__B2 _12337_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13245_ _13320_/A VGND VGND VPWR VPWR _13245_/X sky130_fd_sc_hd__buf_2
XFILLER_182_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ _13197_/A _13173_/X _13176_/C VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__and3_4
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15288__B1 _15183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _25476_/Q VGND VGND VPWR VPWR _12127_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24741__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17984_ _17984_/A _23787_/Q VGND VGND VPWR VPWR _17988_/B sky130_fd_sc_hd__or2_4
XFILLER_96_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19723_ _19722_/Y _19720_/X _19656_/X _19720_/X VGND VGND VPWR VPWR _19723_/X sky130_fd_sc_hd__a2bb2o_4
X_12058_ _17456_/A VGND VGND VPWR VPWR _12059_/A sky130_fd_sc_hd__inv_2
X_16935_ _16935_/A VGND VGND VPWR VPWR _17759_/C sky130_fd_sc_hd__inv_2
XFILLER_237_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12510__A1 _12273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19654_ _19650_/Y _19653_/X _19439_/X _19653_/X VGND VGND VPWR VPWR _19654_/X sky130_fd_sc_hd__a2bb2o_4
X_16866_ _20102_/A VGND VGND VPWR VPWR _16866_/X sky130_fd_sc_hd__buf_2
XFILLER_238_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16788__B1 _16534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18605_ _16603_/Y _18604_/X _16603_/Y _18604_/X VGND VGND VPWR VPWR _18605_/X sky130_fd_sc_hd__a2bb2o_4
X_15817_ _12377_/Y _15811_/X _11783_/X _15811_/X VGND VGND VPWR VPWR _15817_/X sky130_fd_sc_hd__a2bb2o_4
X_19585_ _21828_/B _19580_/X _11957_/X _19580_/X VGND VGND VPWR VPWR _23696_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16797_ _16794_/Y _16792_/X _16796_/X _16792_/X VGND VGND VPWR VPWR _16797_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18536_ _18531_/A _18531_/B _18505_/X _18533_/B VGND VGND VPWR VPWR _18537_/A sky130_fd_sc_hd__a211o_4
X_15748_ HWDATA[16] VGND VGND VPWR VPWR _15748_/X sky130_fd_sc_hd__buf_2
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21533__B1 _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18467_ _18467_/A _18517_/A VGND VGND VPWR VPWR _18486_/C sky130_fd_sc_hd__or2_4
XFILLER_61_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15679_ _21170_/A VGND VGND VPWR VPWR _21874_/A sky130_fd_sc_hd__buf_2
X_17418_ _17396_/X _17410_/X _21008_/B _24341_/Q _17413_/X VGND VGND VPWR VPWR _17418_/X
+ sky130_fd_sc_hd__a32o_4
X_18398_ _16250_/Y _24174_/Q _16250_/Y _24174_/Q VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22493__A _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17349_ _17257_/Y _17347_/A VGND VGND VPWR VPWR _17349_/X sky130_fd_sc_hd__or2_4
XFILLER_174_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23038__B1 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20360_ _20360_/A VGND VGND VPWR VPWR _20360_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23101__B _22968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16712__B1 _16530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19019_ _19019_/A VGND VGND VPWR VPWR _19019_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24829__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20291_ _20278_/Y VGND VGND VPWR VPWR _20291_/X sky130_fd_sc_hd__buf_2
X_22030_ _22025_/X _22029_/X _21499_/X VGND VGND VPWR VPWR _22030_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23210__B1 _12888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23981_ _24003_/CLK _23981_/D HRESETn VGND VGND VPWR VPWR _23981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_229_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_31_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_31_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22932_ _16682_/Y _23177_/B VGND VGND VPWR VPWR _22932_/X sky130_fd_sc_hd__and2_4
XFILLER_189_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22863_ _12801_/Y _22530_/B _22861_/X _12568_/Y _22862_/X VGND VGND VPWR VPWR _22863_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_243_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24602_ _24602_/CLK _24602_/D HRESETn VGND VGND VPWR VPWR _24602_/Q sky130_fd_sc_hd__dfrtp_4
X_21814_ _21676_/A _19955_/Y VGND VGND VPWR VPWR _21815_/C sky130_fd_sc_hd__or2_4
X_22794_ _15800_/A _22792_/X _22503_/X _11802_/A _22793_/X VGND VGND VPWR VPWR _22794_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_231_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24533_ _24532_/CLK _24533_/D HRESETn VGND VGND VPWR VPWR _24533_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21745_ _21744_/X VGND VGND VPWR VPWR _21745_/Y sky130_fd_sc_hd__inv_2
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24464_ _24430_/CLK _24464_/D HRESETn VGND VGND VPWR VPWR _24464_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21676_ _21676_/A _21676_/B VGND VGND VPWR VPWR _21677_/C sky130_fd_sc_hd__or2_4
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23415_ _23560_/CLK _20375_/X VGND VGND VPWR VPWR _23415_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22834__C _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20627_ _20627_/A _20624_/A VGND VGND VPWR VPWR _20627_/Y sky130_fd_sc_hd__nand2_4
XFILLER_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_155_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _25177_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24395_ _24407_/CLK _24395_/D HRESETn VGND VGND VPWR VPWR _24395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23346_ _24482_/Q _22673_/B _23190_/X VGND VGND VPWR VPWR _23346_/X sky130_fd_sc_hd__o21a_4
X_20558_ _14455_/Y _20551_/X _20608_/A _20557_/X VGND VGND VPWR VPWR _20559_/A sky130_fd_sc_hd__a211o_4
XFILLER_164_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13517__B1 _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23277_ _21879_/A _23274_/X _23277_/C VGND VGND VPWR VPWR _23277_/X sky130_fd_sc_hd__and3_4
X_20489_ _20486_/Y _20533_/C _20535_/A VGND VGND VPWR VPWR _24090_/D sky130_fd_sc_hd__a21o_4
XFILLER_138_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23044__A3 _22861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13030_ _13029_/X VGND VGND VPWR VPWR _13031_/B sky130_fd_sc_hd__inv_2
X_25016_ _25011_/CLK _15289_/X HRESETn VGND VGND VPWR VPWR _14984_/A sky130_fd_sc_hd__dfrtp_4
X_22228_ _22228_/A _22226_/X _22228_/C VGND VGND VPWR VPWR _22228_/X sky130_fd_sc_hd__and3_4
XANTENNA__21747__A _21747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22159_ _22159_/A _21103_/A VGND VGND VPWR VPWR _22159_/X sky130_fd_sc_hd__or2_4
XANTENNA__23384__D scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14981_ _25033_/Q VGND VGND VPWR VPWR _15075_/D sky130_fd_sc_hd__inv_2
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22555__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16720_ _16720_/A VGND VGND VPWR VPWR _16720_/Y sky130_fd_sc_hd__inv_2
X_13932_ _13951_/A _13951_/B _13950_/A _13952_/C VGND VGND VPWR VPWR _13932_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22578__A _16703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13863_ _13862_/A _13867_/A _13861_/X _13862_/Y VGND VGND VPWR VPWR _25259_/D sky130_fd_sc_hd__a211o_4
X_16651_ _16651_/A VGND VGND VPWR VPWR _23303_/A sky130_fd_sc_hd__inv_2
XFILLER_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16576__A _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__B _22424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _25386_/Q VGND VGND VPWR VPWR _12815_/A sky130_fd_sc_hd__inv_2
X_15602_ _15614_/A VGND VGND VPWR VPWR _15602_/X sky130_fd_sc_hd__buf_2
X_19370_ _19366_/Y _19369_/X _19326_/X _19369_/X VGND VGND VPWR VPWR _19370_/X sky130_fd_sc_hd__a2bb2o_4
X_13794_ _13779_/X _13793_/X _13481_/X _13793_/X VGND VGND VPWR VPWR _25281_/D sky130_fd_sc_hd__a2bb2o_4
X_16582_ _16581_/Y _16579_/X _16412_/X _16579_/X VGND VGND VPWR VPWR _24540_/D sky130_fd_sc_hd__a2bb2o_4
X_18321_ _18320_/X VGND VGND VPWR VPWR _18321_/Y sky130_fd_sc_hd__inv_2
X_12745_ _25407_/Q _12745_/B VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__or2_4
X_15533_ _15544_/A VGND VGND VPWR VPWR _15533_/X sky130_fd_sc_hd__buf_2
XFILLER_203_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_51_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15464_ _13923_/A _15458_/X _15455_/X _13955_/B _15461_/X VGND VGND VPWR VPWR _24968_/D
+ sky130_fd_sc_hd__a32o_4
X_18252_ _18243_/A VGND VGND VPWR VPWR _18252_/X sky130_fd_sc_hd__buf_2
XANTENNA__23268__B1 _16925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12676_ _12596_/Y _12676_/B VGND VGND VPWR VPWR _12676_/X sky130_fd_sc_hd__or2_4
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16942__B1 _16143_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14415_/A _14388_/B VGND VGND VPWR VPWR _14415_/X sky130_fd_sc_hd__or2_4
X_17203_ _24375_/Q VGND VGND VPWR VPWR _17203_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _15394_/X VGND VGND VPWR VPWR _24993_/D sky130_fd_sc_hd__inv_2
X_18183_ _14656_/A _18181_/X _18183_/C VGND VGND VPWR VPWR _18183_/X sky130_fd_sc_hd__and3_4
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _25169_/Q VGND VGND VPWR VPWR _14349_/A sky130_fd_sc_hd__inv_2
X_17134_ _17129_/A _17129_/B _17130_/Y _17065_/X VGND VGND VPWR VPWR _17135_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13508__B1 _11834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17065_ _17393_/B VGND VGND VPWR VPWR _17065_/X sky130_fd_sc_hd__buf_2
XANTENNA__24922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14277_ _14277_/A VGND VGND VPWR VPWR _14277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11791__A1_N _11789_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22760__B _22610_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16016_ _24748_/Q VGND VGND VPWR VPWR _16016_/Y sky130_fd_sc_hd__inv_2
X_13228_ _13228_/A VGND VGND VPWR VPWR _13385_/A sky130_fd_sc_hd__buf_2
XANTENNA__20254__B1 _19761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13159_ _13212_/A VGND VGND VPWR VPWR _13271_/A sky130_fd_sc_hd__inv_2
XFILLER_112_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17967_ _17941_/A _17965_/X _17967_/C VGND VGND VPWR VPWR _17967_/X sky130_fd_sc_hd__and3_4
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19706_ _13326_/B VGND VGND VPWR VPWR _19706_/Y sky130_fd_sc_hd__inv_2
X_16918_ _24287_/Q VGND VGND VPWR VPWR _17753_/B sky130_fd_sc_hd__inv_2
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17898_ _17710_/X _17898_/B VGND VGND VPWR VPWR _17899_/A sky130_fd_sc_hd__and2_4
XFILLER_238_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19637_ _19635_/Y _19633_/X _19636_/X _19633_/X VGND VGND VPWR VPWR _19637_/X sky130_fd_sc_hd__a2bb2o_4
X_16849_ _16853_/A VGND VGND VPWR VPWR _16849_/X sky130_fd_sc_hd__buf_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15433__B1 _15324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19568_ _19568_/A VGND VGND VPWR VPWR _19568_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12798__A1 _25375_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18519_ _18467_/A _18517_/X _18518_/Y VGND VGND VPWR VPWR _18519_/X sky130_fd_sc_hd__o21a_4
XFILLER_34_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19797__A _19788_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19499_ _21501_/B _19496_/X _11964_/X _19496_/X VGND VGND VPWR VPWR _19499_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21530_ _22721_/B VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__buf_2
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23112__A _23089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21461_ _22810_/A _21439_/Y _21454_/Y _21455_/X _21460_/X VGND VGND VPWR VPWR _21461_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_228_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _25253_/CLK sky130_fd_sc_hd__clkbuf_1
X_23200_ _23052_/X _23199_/X _22986_/X _12536_/A _23120_/X VGND VGND VPWR VPWR _23201_/B
+ sky130_fd_sc_hd__a32o_4
X_20412_ _20410_/Y _20411_/Y _11851_/A _20411_/Y VGND VGND VPWR VPWR _23401_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17489__A1 _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24180_ _24523_/CLK _24180_/D HRESETn VGND VGND VPWR VPWR _24180_/Q sky130_fd_sc_hd__dfrtp_4
X_21392_ _14687_/A _21392_/B _21391_/X VGND VGND VPWR VPWR _21392_/X sky130_fd_sc_hd__and3_4
X_23131_ _23123_/X _23127_/Y _22881_/X _23130_/X VGND VGND VPWR VPWR _23131_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24663__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20343_ _21380_/A VGND VGND VPWR VPWR _20343_/X sky130_fd_sc_hd__buf_2
XANTENNA__23241__A2_N _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23062_ _22986_/A VGND VGND VPWR VPWR _23062_/X sky130_fd_sc_hd__buf_2
XFILLER_150_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20274_ _13446_/B VGND VGND VPWR VPWR _20274_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22013_ _21972_/B VGND VGND VPWR VPWR _22013_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15565__A _21855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23195__C1 _23194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23964_ _23946_/CLK _23964_/D HRESETn VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22915_ _23056_/A _22914_/X VGND VGND VPWR VPWR _22923_/C sky130_fd_sc_hd__and2_4
XFILLER_244_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23895_ _24101_/CLK _23895_/D VGND VGND VPWR VPWR _19019_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22846_ _16687_/Y _22808_/A _15604_/Y _22845_/X VGND VGND VPWR VPWR _22846_/X sky130_fd_sc_hd__o22a_4
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12789__A1 _25392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22777_ _21126_/B VGND VGND VPWR VPWR _22777_/X sky130_fd_sc_hd__buf_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22170__B1 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12529_/Y VGND VGND VPWR VPWR _12618_/B sky130_fd_sc_hd__buf_2
X_24516_ _24684_/CLK _24516_/D HRESETn VGND VGND VPWR VPWR _24516_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_38_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21728_ _14432_/Y _14232_/A _14455_/Y _15471_/A VGND VGND VPWR VPWR _21730_/C sky130_fd_sc_hd__o22a_4
XFILLER_212_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25496_ _24171_/CLK _12048_/X HRESETn VGND VGND VPWR VPWR _12047_/A sky130_fd_sc_hd__dfrtp_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12461_ _12247_/X _12440_/C VGND VGND VPWR VPWR _12464_/B sky130_fd_sc_hd__or2_4
X_24447_ _25043_/CLK _16813_/X HRESETn VGND VGND VPWR VPWR _14976_/A sky130_fd_sc_hd__dfrtp_4
X_21659_ _22549_/B _21658_/X _13574_/Y _22549_/B VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14200_ _11731_/A _19594_/B _11734_/B _13786_/A VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__or4_4
XFILLER_200_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18116__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15180_ _15067_/A _15172_/X VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__and2_4
XFILLER_137_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12392_ _12391_/X VGND VGND VPWR VPWR _13017_/B sky130_fd_sc_hd__buf_2
X_24378_ _24378_/CLK _24378_/D HRESETn VGND VGND VPWR VPWR _24378_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22861__A _21719_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14131_ _23968_/Q VGND VGND VPWR VPWR _14131_/X sky130_fd_sc_hd__buf_2
XFILLER_138_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23329_ _22563_/X _23328_/X _22145_/C _25556_/Q _22565_/X VGND VGND VPWR VPWR _23329_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_193_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17955__A _18023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _14062_/A _14056_/Y _14062_/C VGND VGND VPWR VPWR _14063_/A sky130_fd_sc_hd__or3_4
XFILLER_153_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _25371_/Q _13013_/B VGND VGND VPWR VPWR _13015_/B sky130_fd_sc_hd__or2_4
XANTENNA__20236__B1 _19817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18870_ _16482_/A _18702_/A _24572_/Q _18696_/D VGND VGND VPWR VPWR _18871_/D sky130_fd_sc_hd__a2bb2o_4
X_17821_ _16950_/Y _17820_/X VGND VGND VPWR VPWR _17824_/B sky130_fd_sc_hd__or2_4
XFILLER_95_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24003__D sda_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17752_ _17752_/A VGND VGND VPWR VPWR _17753_/A sky130_fd_sc_hd__inv_2
X_14964_ _14964_/A VGND VGND VPWR VPWR _14965_/A sky130_fd_sc_hd__inv_2
X_16703_ _24494_/Q VGND VGND VPWR VPWR _16703_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13915_ _13915_/A _13955_/B _13963_/A _13911_/Y VGND VGND VPWR VPWR _13916_/A sky130_fd_sc_hd__or4_4
XFILLER_35_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17683_ _17687_/A _17683_/B _17682_/Y VGND VGND VPWR VPWR _24306_/D sky130_fd_sc_hd__and3_4
X_14895_ _15070_/A VGND VGND VPWR VPWR _14895_/X sky130_fd_sc_hd__buf_2
XANTENNA__25192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19422_ _19415_/A VGND VGND VPWR VPWR _19422_/X sky130_fd_sc_hd__buf_2
X_16634_ _16633_/X VGND VGND VPWR VPWR _16634_/Y sky130_fd_sc_hd__inv_2
X_13846_ _11847_/A VGND VGND VPWR VPWR _13846_/X sky130_fd_sc_hd__buf_2
XFILLER_235_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19353_ _19353_/A VGND VGND VPWR VPWR _19353_/X sky130_fd_sc_hd__buf_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13777_ _13757_/A _14712_/A _13775_/X VGND VGND VPWR VPWR _13777_/X sky130_fd_sc_hd__o21a_4
X_16565_ _16564_/Y _16560_/X _16395_/X _16560_/X VGND VGND VPWR VPWR _24547_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18304_ _21509_/A _18303_/X _21509_/A _18303_/X VGND VGND VPWR VPWR _24220_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22755__B _21104_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15516_ _15515_/Y _15513_/X HADDR[16] _15513_/X VGND VGND VPWR VPWR _15516_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19410__A _19139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12728_ _12728_/A _12715_/X _12727_/Y VGND VGND VPWR VPWR _25413_/D sky130_fd_sc_hd__and3_4
X_19284_ _19283_/Y _19281_/X _16876_/X _19281_/X VGND VGND VPWR VPWR _19284_/X sky130_fd_sc_hd__a2bb2o_4
X_16496_ _16494_/Y _16495_/X _16410_/X _16495_/X VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18235_ _18107_/A _18227_/X _18235_/C VGND VGND VPWR VPWR _18235_/X sky130_fd_sc_hd__and3_4
XFILLER_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12659_ _12710_/B _12627_/X _12588_/Y _12628_/A VGND VGND VPWR VPWR _12660_/B sky130_fd_sc_hd__or4_4
X_15447_ _15447_/A VGND VGND VPWR VPWR _15447_/X sky130_fd_sc_hd__buf_2
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18166_ _18166_/A _18166_/B _18166_/C VGND VGND VPWR VPWR _18170_/B sky130_fd_sc_hd__and3_4
XFILLER_156_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18668__B1 _24521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15378_ _15306_/B _15381_/B VGND VGND VPWR VPWR _15378_/Y sky130_fd_sc_hd__nand2_4
XFILLER_156_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22771__A _21890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17117_ _17106_/A _17117_/B _17117_/C VGND VGND VPWR VPWR _24396_/D sky130_fd_sc_hd__and3_4
X_14329_ _14315_/A _14328_/X _13497_/A _14320_/X VGND VGND VPWR VPWR _25178_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18097_ _18097_/A VGND VGND VPWR VPWR _18166_/A sky130_fd_sc_hd__buf_2
XFILLER_171_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_58_0_HCLK clkbuf_8_58_0_HCLK/A VGND VGND VPWR VPWR _24230_/CLK sky130_fd_sc_hd__clkbuf_1
X_17048_ _24381_/Q VGND VGND VPWR VPWR _17048_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24958__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18999_ _19139_/A VGND VGND VPWR VPWR _18999_/X sky130_fd_sc_hd__buf_2
XFILLER_86_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21834__B _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19640__A1_N _19638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20961_ _13676_/A _20956_/A _20952_/A VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__or3_4
XFILLER_39_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22011__A _13793_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22700_ _20756_/Y _23144_/A _15611_/Y _22289_/X VGND VGND VPWR VPWR _22700_/X sky130_fd_sc_hd__o22a_4
X_23680_ _23799_/CLK _19640_/X VGND VGND VPWR VPWR _19638_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_226_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _13672_/A _13671_/X VGND VGND VPWR VPWR _20896_/A sky130_fd_sc_hd__or2_4
XFILLER_242_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22631_ _22631_/A _22468_/X VGND VGND VPWR VPWR _22631_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22152__B1 _22810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22665__B _22662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25350_ _25368_/CLK _25350_/D HRESETn VGND VGND VPWR VPWR _25350_/Q sky130_fd_sc_hd__dfrtp_4
X_22562_ _15715_/X VGND VGND VPWR VPWR _22562_/X sky130_fd_sc_hd__buf_2
XFILLER_194_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24301_ _23590_/CLK _24301_/D HRESETn VGND VGND VPWR VPWR _17538_/A sky130_fd_sc_hd__dfrtp_4
X_21513_ _13826_/X VGND VGND VPWR VPWR _21513_/X sky130_fd_sc_hd__buf_2
XFILLER_210_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24844__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25281_ _25281_/CLK _25281_/D HRESETn VGND VGND VPWR VPWR _13778_/A sky130_fd_sc_hd__dfrtp_4
X_22493_ _22437_/X VGND VGND VPWR VPWR _22493_/X sky130_fd_sc_hd__buf_2
X_24232_ _24238_/CLK _24232_/D HRESETn VGND VGND VPWR VPWR _24232_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21444_ _21444_/A _23016_/A VGND VGND VPWR VPWR _21444_/X sky130_fd_sc_hd__or2_4
XFILLER_166_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24163_ _24192_/CLK _18603_/Y HRESETn VGND VGND VPWR VPWR _24163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17775__A _16925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21375_ _21375_/A VGND VGND VPWR VPWR _21375_/X sky130_fd_sc_hd__buf_2
X_23114_ _24778_/Q _23158_/B VGND VGND VPWR VPWR _23114_/X sky130_fd_sc_hd__or2_4
XFILLER_162_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20326_ _20326_/A VGND VGND VPWR VPWR _22253_/B sky130_fd_sc_hd__inv_2
XFILLER_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21297__A _21877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24094_ _24095_/CLK _24094_/D HRESETn VGND VGND VPWR VPWR _20445_/A sky130_fd_sc_hd__dfstp_4
XFILLER_162_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15893__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23045_ _22771_/X _23043_/X _22702_/X _23044_/X VGND VGND VPWR VPWR _23045_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20257_ _20256_/X VGND VGND VPWR VPWR _20270_/A sky130_fd_sc_hd__inv_2
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20188_ _20188_/A VGND VGND VPWR VPWR _20188_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24996_ _24981_/CLK _24996_/D HRESETn VGND VGND VPWR VPWR _15383_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11961_ _19643_/A VGND VGND VPWR VPWR _11961_/X sky130_fd_sc_hd__buf_2
XFILLER_245_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15660__A3 _15656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23947_ _23395_/CLK _20995_/B HRESETn VGND VGND VPWR VPWR _20419_/B sky130_fd_sc_hd__dfstp_4
XFILLER_57_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ _11666_/Y _13700_/B VGND VGND VPWR VPWR _13707_/B sky130_fd_sc_hd__or2_4
XFILLER_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20206__A2_N _20205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14680_ _19436_/B VGND VGND VPWR VPWR _19166_/B sky130_fd_sc_hd__buf_2
XFILLER_245_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11892_ _11887_/A VGND VGND VPWR VPWR _11892_/Y sky130_fd_sc_hd__inv_2
X_23878_ _23459_/CLK _23878_/D VGND VGND VPWR VPWR _23878_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_232_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18864__A1_N _16512_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22856__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _13625_/X _13630_/X _13625_/X _13630_/X VGND VGND VPWR VPWR _14801_/B sky130_fd_sc_hd__a2bb2o_4
X_22829_ _22684_/B VGND VGND VPWR VPWR _22830_/C sky130_fd_sc_hd__buf_2
XFILLER_204_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13562_ _13560_/Y _25094_/Q _25261_/Q _13561_/Y VGND VGND VPWR VPWR _13563_/D sky130_fd_sc_hd__a2bb2o_4
X_16350_ _16348_/Y _16346_/X _16349_/X _16346_/X VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__a2bb2o_4
X_25548_ _24697_/CLK _25548_/D HRESETn VGND VGND VPWR VPWR _25548_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12513_ _12513_/A _12478_/B VGND VGND VPWR VPWR _12513_/Y sky130_fd_sc_hd__nand2_4
X_15301_ _15388_/A VGND VGND VPWR VPWR _15337_/A sky130_fd_sc_hd__buf_2
X_16281_ _15655_/X _16288_/B _16090_/X _21021_/A _16280_/X VGND VGND VPWR VPWR _24651_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_40_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24585__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ _13493_/A VGND VGND VPWR VPWR _13493_/Y sky130_fd_sc_hd__inv_2
X_25479_ _24196_/CLK _25479_/D HRESETn VGND VGND VPWR VPWR _25479_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18020_ _18013_/A VGND VGND VPWR VPWR _18129_/A sky130_fd_sc_hd__buf_2
XFILLER_185_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12444_ _12293_/A _12444_/B VGND VGND VPWR VPWR _12444_/X sky130_fd_sc_hd__or2_4
X_15232_ _15232_/A _15231_/X VGND VGND VPWR VPWR _15232_/X sky130_fd_sc_hd__or2_4
XFILLER_200_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_211_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24601_/CLK sky130_fd_sc_hd__clkbuf_1
X_15163_ _15162_/Y _24588_/Q _15311_/A _15134_/Y VGND VGND VPWR VPWR _15170_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _24845_/Q VGND VGND VPWR VPWR _12375_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14114_ _25230_/Q VGND VGND VPWR VPWR _14114_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15094_ _15380_/A _24601_/Q _15092_/Y _24601_/Q VGND VGND VPWR VPWR _15103_/A sky130_fd_sc_hd__a2bb2o_4
X_19971_ _19971_/A VGND VGND VPWR VPWR _22034_/B sky130_fd_sc_hd__inv_2
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15884__B1 _11776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14045_ _23941_/Q _14040_/Y _14045_/C VGND VGND VPWR VPWR _14060_/B sky130_fd_sc_hd__or3_4
X_18922_ _18916_/Y VGND VGND VPWR VPWR _18922_/X sky130_fd_sc_hd__buf_2
X_18853_ _16504_/Y _18768_/A _24573_/Q _18756_/A VGND VGND VPWR VPWR _18856_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18822__B1 _18714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17804_ _17753_/B _17803_/X VGND VGND VPWR VPWR _17807_/B sky130_fd_sc_hd__or2_4
XFILLER_79_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15933__A _19761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18784_ _18776_/A _18784_/B _18784_/C VGND VGND VPWR VPWR _24144_/D sky130_fd_sc_hd__and3_4
X_15996_ _12233_/Y _15990_/X _15995_/X _15990_/X VGND VGND VPWR VPWR _24755_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17735_ _17733_/A _17720_/X _17734_/Y VGND VGND VPWR VPWR _17735_/X sky130_fd_sc_hd__o21a_4
XFILLER_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14947_ _25015_/Q _24421_/Q _15290_/A _14946_/Y VGND VGND VPWR VPWR _14947_/X sky130_fd_sc_hd__o22a_4
XFILLER_224_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17666_ _17666_/A _17666_/B VGND VGND VPWR VPWR _17666_/X sky130_fd_sc_hd__or2_4
X_14878_ _14873_/A VGND VGND VPWR VPWR _14878_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22766__A _16691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19391_/X VGND VGND VPWR VPWR _19405_/X sky130_fd_sc_hd__buf_2
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16617_ _16617_/A VGND VGND VPWR VPWR _16617_/Y sky130_fd_sc_hd__inv_2
X_13829_ _13828_/X VGND VGND VPWR VPWR _13848_/A sky130_fd_sc_hd__buf_2
X_17597_ _17596_/A _17596_/B VGND VGND VPWR VPWR _17597_/Y sky130_fd_sc_hd__nand2_4
XFILLER_90_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19336_ _19335_/Y _19331_/X _19246_/X _19331_/X VGND VGND VPWR VPWR _23784_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16548_ _24552_/Q VGND VGND VPWR VPWR _16548_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22685__A1 _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_21_0_HCLK clkbuf_5_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19267_ _21896_/B _19264_/X _16885_/X _19264_/X VGND VGND VPWR VPWR _23809_/D sky130_fd_sc_hd__a2bb2o_4
X_16479_ _16478_/Y _16476_/X _16393_/X _16476_/X VGND VGND VPWR VPWR _16479_/X sky130_fd_sc_hd__a2bb2o_4
X_18218_ _17975_/X _18216_/X _18217_/X VGND VGND VPWR VPWR _18218_/X sky130_fd_sc_hd__and3_4
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19198_ _23833_/Q VGND VGND VPWR VPWR _19198_/Y sky130_fd_sc_hd__inv_2
X_18149_ _17977_/A _18149_/B VGND VGND VPWR VPWR _18149_/X sky130_fd_sc_hd__or2_4
XFILLER_191_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21829__B _19638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21160_ _21160_/A VGND VGND VPWR VPWR _21160_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12809__A2_N _22641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20111_ _23513_/Q VGND VGND VPWR VPWR _21925_/B sky130_fd_sc_hd__inv_2
XFILLER_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19066__B1 _18991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21091_ _21091_/A _21091_/B VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__or2_4
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20042_ _22271_/B _20039_/X _19993_/X _20039_/X VGND VGND VPWR VPWR _23539_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21845__A _22947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15627__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24850_ _24878_/CLK _24850_/D HRESETn VGND VGND VPWR VPWR _24850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23801_ _23577_/CLK _23801_/D VGND VGND VPWR VPWR _23801_/Q sky130_fd_sc_hd__dfxtp_4
X_24781_ _24781_/CLK _15951_/X HRESETn VGND VGND VPWR VPWR _23228_/A sky130_fd_sc_hd__dfrtp_4
X_21993_ _21990_/X _21991_/X _21992_/X VGND VGND VPWR VPWR _21993_/Y sky130_fd_sc_hd__o21ai_4
XPHY_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23732_ _23555_/CLK _19485_/X VGND VGND VPWR VPWR _19479_/A sky130_fd_sc_hd__dfxtp_4
X_20944_ _20944_/A _20944_/B _13674_/X VGND VGND VPWR VPWR _20949_/B sky130_fd_sc_hd__or3_4
XPHY_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16052__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_207_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23654_/CLK _23663_/D VGND VGND VPWR VPWR _13393_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ _20874_/Y _20870_/X _13668_/X VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__o21a_4
XFILLER_241_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _22562_/X _22613_/X _22144_/A _11824_/A _22940_/A VGND VGND VPWR VPWR _22614_/X
+ sky130_fd_sc_hd__a32o_4
X_25402_ _25402_/CLK _25402_/D HRESETn VGND VGND VPWR VPWR _12790_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23560_/CLK _23594_/D VGND VGND VPWR VPWR _19887_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_241_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25333_ _25488_/CLK _13409_/X HRESETn VGND VGND VPWR VPWR _25333_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22140__A3 _21550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22545_ _22544_/X VGND VGND VPWR VPWR _22545_/X sky130_fd_sc_hd__buf_2
XFILLER_139_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25264_ _25309_/CLK _25264_/D HRESETn VGND VGND VPWR VPWR _25264_/Q sky130_fd_sc_hd__dfrtp_4
X_22476_ _22476_/A _22476_/B VGND VGND VPWR VPWR _22480_/C sky130_fd_sc_hd__nor2_4
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16605__A1_N _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24215_ _23522_/CLK _18338_/Y HRESETn VGND VGND VPWR VPWR _17464_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21427_ _21427_/A VGND VGND VPWR VPWR _22810_/A sky130_fd_sc_hd__buf_2
X_25195_ _25200_/CLK _14274_/X HRESETn VGND VGND VPWR VPWR _14272_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21100__A1 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12160_ _12160_/A _12157_/A VGND VGND VPWR VPWR _12162_/A sky130_fd_sc_hd__and2_4
X_24146_ _24966_/CLK _24146_/D HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21358_ _21357_/X VGND VGND VPWR VPWR _21358_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_41_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23514_/CLK sky130_fd_sc_hd__clkbuf_1
X_20309_ _20307_/Y _20303_/X _19996_/X _20308_/X VGND VGND VPWR VPWR _23441_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12091_ _12090_/Y _12088_/X _11856_/X _12088_/X VGND VGND VPWR VPWR _12091_/X sky130_fd_sc_hd__a2bb2o_4
X_24077_ _24073_/CLK _24077_/D HRESETn VGND VGND VPWR VPWR _20964_/A sky130_fd_sc_hd__dfrtp_4
X_21289_ _21279_/X _21286_/X _21288_/X VGND VGND VPWR VPWR _21290_/D sky130_fd_sc_hd__a21o_4
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23028_ _16028_/A _21039_/X _21068_/X _23027_/X VGND VGND VPWR VPWR _23029_/C sky130_fd_sc_hd__a211o_4
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15850_ _15833_/X _15844_/X _15782_/X _24825_/Q _15802_/A VGND VGND VPWR VPWR _24825_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18280__A1 _13793_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15094__B2 _24601_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14801_ _14801_/A _14801_/B _14801_/C _14801_/D VGND VGND VPWR VPWR _14801_/X sky130_fd_sc_hd__or4_4
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15781_ HWDATA[0] VGND VGND VPWR VPWR _19761_/A sky130_fd_sc_hd__buf_2
X_12993_ _12992_/Y VGND VGND VPWR VPWR _13021_/C sky130_fd_sc_hd__buf_2
X_24979_ _24979_/CLK _15448_/X HRESETn VGND VGND VPWR VPWR _24979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17520_ _24320_/Q VGND VGND VPWR VPWR _17520_/Y sky130_fd_sc_hd__inv_2
X_14732_ _14731_/X VGND VGND VPWR VPWR _14732_/Y sky130_fd_sc_hd__inv_2
X_11944_ _11934_/X VGND VGND VPWR VPWR _11944_/X sky130_fd_sc_hd__buf_2
XFILLER_206_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21490__A _21687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17451_ _13818_/A VGND VGND VPWR VPWR _19139_/A sky130_fd_sc_hd__buf_2
XANTENNA__24766__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ _13818_/A VGND VGND VPWR VPWR _13481_/A sky130_fd_sc_hd__buf_2
X_14663_ _13614_/B _14650_/C _17945_/A _14662_/X VGND VGND VPWR VPWR _25081_/D sky130_fd_sc_hd__a22oi_4
XFILLER_221_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16402_ HWDATA[24] VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__buf_2
X_13614_ _14794_/A _13614_/B VGND VGND VPWR VPWR _13615_/A sky130_fd_sc_hd__and2_4
X_17382_ _17363_/A _17378_/B _17381_/X VGND VGND VPWR VPWR _24351_/D sky130_fd_sc_hd__and3_4
X_14594_ _14590_/B _14566_/X _14593_/X _13779_/X _14593_/A VGND VGND VPWR VPWR _25100_/D
+ sky130_fd_sc_hd__a32o_4
X_19121_ _19134_/A VGND VGND VPWR VPWR _19121_/X sky130_fd_sc_hd__buf_2
XFILLER_41_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16333_ _16352_/A VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__buf_2
X_13545_ _25308_/Q VGND VGND VPWR VPWR _13652_/A sky130_fd_sc_hd__inv_2
XANTENNA__16734__D _21173_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19052_ _23884_/Q VGND VGND VPWR VPWR _19052_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13476_ _12059_/A _16378_/B _15791_/C _13476_/D VGND VGND VPWR VPWR _21577_/B sky130_fd_sc_hd__or4_4
X_16264_ _16264_/A VGND VGND VPWR VPWR _16264_/X sky130_fd_sc_hd__buf_2
XFILLER_186_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18003_ _18234_/A _17996_/X _18003_/C VGND VGND VPWR VPWR _18004_/C sky130_fd_sc_hd__or3_4
X_12427_ _25463_/Q _12427_/B VGND VGND VPWR VPWR _12429_/B sky130_fd_sc_hd__or2_4
X_15215_ _14996_/A _15215_/B _15215_/C VGND VGND VPWR VPWR _15215_/X sky130_fd_sc_hd__or3_4
XFILLER_145_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16195_ _16382_/A _16468_/B VGND VGND VPWR VPWR _16202_/A sky130_fd_sc_hd__nor2_4
X_12358_ _12358_/A VGND VGND VPWR VPWR _12997_/D sky130_fd_sc_hd__inv_2
X_15146_ _24998_/Q VGND VGND VPWR VPWR _15306_/B sky130_fd_sc_hd__inv_2
XANTENNA__25554__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15077_ _14962_/A _14956_/Y _15075_/X _15077_/D VGND VGND VPWR VPWR _15078_/B sky130_fd_sc_hd__or4_4
X_19954_ _19953_/Y _19951_/X _19636_/X _19951_/X VGND VGND VPWR VPWR _23569_/D sky130_fd_sc_hd__a2bb2o_4
X_12289_ _25439_/Q VGND VGND VPWR VPWR _12513_/A sky130_fd_sc_hd__inv_2
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14028_ _14028_/A _14027_/D _14027_/A _14028_/D VGND VGND VPWR VPWR _14028_/X sky130_fd_sc_hd__or4_4
X_18905_ _20079_/A _20079_/B _20079_/C _18905_/D VGND VGND VPWR VPWR _18905_/X sky130_fd_sc_hd__or4_4
X_19885_ _23595_/Q VGND VGND VPWR VPWR _19885_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18836_ _16485_/Y _18737_/A _16485_/Y _18737_/A VGND VGND VPWR VPWR _18840_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11894__A1 _11890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18767_ _18764_/B VGND VGND VPWR VPWR _18768_/B sky130_fd_sc_hd__inv_2
X_15979_ _15974_/X _15977_/X _16241_/A _24767_/Q _15975_/X VGND VGND VPWR VPWR _15979_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21659__A1_N _22549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17718_ _17717_/X VGND VGND VPWR VPWR _18289_/A sky130_fd_sc_hd__inv_2
X_18698_ _18765_/A _18764_/A _18698_/C _18763_/A VGND VGND VPWR VPWR _18752_/A sky130_fd_sc_hd__or4_4
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16034__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22496__A _24626_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17649_ _17646_/C _17646_/D VGND VGND VPWR VPWR _17649_/X sky130_fd_sc_hd__or2_4
XFILLER_223_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16494__A _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _17404_/A _17404_/B VGND VGND VPWR VPWR _20660_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22658__A1 _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19319_ _19318_/Y _19316_/X _19184_/X _19316_/X VGND VGND VPWR VPWR _19319_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20591_ _20591_/A VGND VGND VPWR VPWR _20591_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22330_ _11999_/Y _12106_/A _11998_/Y _12080_/A VGND VGND VPWR VPWR _22330_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23120__A _21436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22261_ _22264_/A _20019_/Y VGND VGND VPWR VPWR _22261_/X sky130_fd_sc_hd__or2_4
X_24000_ _24000_/CLK _20680_/Y HRESETn VGND VGND VPWR VPWR _24000_/Q sky130_fd_sc_hd__dfrtp_4
X_21212_ _21212_/A _21212_/B _21212_/C VGND VGND VPWR VPWR _21212_/X sky130_fd_sc_hd__and3_4
XFILLER_247_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22192_ _22192_/A VGND VGND VPWR VPWR _22192_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_0_0_HCLK clkbuf_7_0_0_HCLK/X VGND VGND VPWR VPWR _23716_/CLK sky130_fd_sc_hd__clkbuf_1
X_21143_ _21143_/A _21138_/X _21141_/X _21143_/D VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__and4_4
XFILLER_144_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_28_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21074_ _21747_/A _21073_/Y _24718_/Q _21747_/A VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20025_ _21944_/B _20022_/X _20000_/X _20022_/X VGND VGND VPWR VPWR _23545_/D sky130_fd_sc_hd__a2bb2o_4
X_24902_ _24020_/CLK _24902_/D HRESETn VGND VGND VPWR VPWR _24902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_219_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24833_ _24849_/CLK _24833_/D HRESETn VGND VGND VPWR VPWR _12327_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24101__D _20969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _14624_/A _21976_/B VGND VGND VPWR VPWR _21976_/X sky130_fd_sc_hd__and2_4
X_24764_ _24756_/CLK _24764_/D HRESETn VGND VGND VPWR VPWR _22608_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16025__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _20836_/A VGND VGND VPWR VPWR _20927_/X sky130_fd_sc_hd__buf_2
X_23715_ _23716_/CLK _23715_/D VGND VGND VPWR VPWR _23715_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19762__B2 _19742_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24695_ _24689_/CLK _24695_/D HRESETn VGND VGND VPWR VPWR _22502_/A sky130_fd_sc_hd__dfrtp_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11660_/A VGND VGND VPWR VPWR _11979_/C sky130_fd_sc_hd__buf_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _20858_/A VGND VGND VPWR VPWR _20858_/Y sky130_fd_sc_hd__inv_2
X_23646_ _23647_/CLK _23646_/D VGND VGND VPWR VPWR _13432_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23577_ _23577_/CLK _19934_/X VGND VGND VPWR VPWR _23577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_179_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20789_ _20789_/A VGND VGND VPWR VPWR _20789_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13290_/X _13330_/B _13329_/X VGND VGND VPWR VPWR _13331_/C sky130_fd_sc_hd__and3_4
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _22527_/X VGND VGND VPWR VPWR _22528_/X sky130_fd_sc_hd__buf_2
X_25316_ _25316_/CLK _25316_/D HRESETn VGND VGND VPWR VPWR _12009_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13443_/A VGND VGND VPWR VPWR _13372_/A sky130_fd_sc_hd__buf_2
XANTENNA__15748__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _22459_/A VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__buf_2
X_25247_ _25246_/CLK _25247_/D HRESETn VGND VGND VPWR VPWR _25247_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14652__A _14650_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12212_ _12212_/A VGND VGND VPWR VPWR _12212_/X sky130_fd_sc_hd__buf_2
X_15000_ _24456_/Q VGND VGND VPWR VPWR _15000_/Y sky130_fd_sc_hd__inv_2
X_13192_ _13192_/A _20255_/A VGND VGND VPWR VPWR _13193_/C sky130_fd_sc_hd__or2_4
X_25178_ _25181_/CLK _25178_/D HRESETn VGND VGND VPWR VPWR _25178_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22821__A1 _16506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15839__B1 _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12143_ _12142_/X VGND VGND VPWR VPWR _12143_/Y sky130_fd_sc_hd__inv_2
X_24129_ _23946_/CLK _24129_/D HRESETn VGND VGND VPWR VPWR _24129_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_151_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21485__A _21485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12074_ _13821_/B VGND VGND VPWR VPWR _21577_/A sky130_fd_sc_hd__buf_2
X_16951_ _16110_/Y _24289_/Q _24706_/Q _16950_/Y VGND VGND VPWR VPWR _16954_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21388__A1 _13547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15902_ _15863_/X VGND VGND VPWR VPWR _15902_/X sky130_fd_sc_hd__buf_2
XFILLER_238_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15483__A _14412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19670_ _19669_/Y _19667_/X _19454_/X _19667_/X VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16882_ _16880_/Y _16877_/X _16881_/X _16877_/X VGND VGND VPWR VPWR _16882_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18621_ _18686_/A VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__buf_2
X_15833_ _22891_/B VGND VGND VPWR VPWR _15833_/X sky130_fd_sc_hd__buf_2
XANTENNA__24947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22337__B1 _20681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18552_ _24178_/Q _18552_/B VGND VGND VPWR VPWR _18552_/X sky130_fd_sc_hd__or2_4
X_15764_ _12532_/Y _15763_/X _11831_/X _15763_/X VGND VGND VPWR VPWR _24870_/D sky130_fd_sc_hd__a2bb2o_4
X_12976_ _12984_/A _12969_/B _12975_/X VGND VGND VPWR VPWR _25378_/D sky130_fd_sc_hd__and3_4
XFILLER_218_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17503_ _11715_/Y _17596_/A _11715_/Y _17596_/A VGND VGND VPWR VPWR _17503_/X sky130_fd_sc_hd__a2bb2o_4
X_14715_ _14714_/X VGND VGND VPWR VPWR _14715_/X sky130_fd_sc_hd__buf_2
XFILLER_205_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11927_ _11885_/A _11929_/A _11919_/X _11926_/Y VGND VGND VPWR VPWR _25517_/D sky130_fd_sc_hd__o22a_4
X_18483_ _18476_/X _18479_/X _18482_/X VGND VGND VPWR VPWR _18557_/B sky130_fd_sc_hd__or3_4
XFILLER_206_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15695_ _13548_/A _15692_/Y _15694_/X _13601_/B VGND VGND VPWR VPWR _15696_/C sky130_fd_sc_hd__a211o_4
X_17434_ _17426_/A VGND VGND VPWR VPWR _17434_/X sky130_fd_sc_hd__buf_2
X_14646_ _13625_/X VGND VGND VPWR VPWR _17941_/A sky130_fd_sc_hd__buf_2
X_11858_ _11853_/Y _11845_/X _11856_/X _11857_/X VGND VGND VPWR VPWR _25529_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17365_ _17359_/C _17364_/X _17298_/A _17361_/B VGND VGND VPWR VPWR _17366_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16464__D _21173_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11789_ _25545_/Q VGND VGND VPWR VPWR _11789_/Y sky130_fd_sc_hd__inv_2
X_14577_ _14601_/A _14577_/B VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__or2_4
XFILLER_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19104_ _23866_/Q VGND VGND VPWR VPWR _22078_/B sky130_fd_sc_hd__inv_2
XANTENNA__22763__B _23053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16316_ _16314_/Y _16312_/X _16315_/X _16312_/X VGND VGND VPWR VPWR _24640_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13528_ _14299_/B VGND VGND VPWR VPWR _13529_/A sky130_fd_sc_hd__buf_2
X_17296_ _17296_/A VGND VGND VPWR VPWR _17298_/A sky130_fd_sc_hd__buf_2
XANTENNA__17857__B _17562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20564__A _14116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19035_ _19034_/Y _19030_/X _19008_/X _19030_/X VGND VGND VPWR VPWR _23891_/D sky130_fd_sc_hd__a2bb2o_4
X_16247_ _24664_/Q VGND VGND VPWR VPWR _16247_/Y sky130_fd_sc_hd__inv_2
X_13459_ _13322_/A _13459_/B _13458_/X VGND VGND VPWR VPWR _13459_/X sky130_fd_sc_hd__and3_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14562__A HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21076__B1 _21882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20418__A3 _13481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16178_ _14779_/A _14769_/X VGND VGND VPWR VPWR _16179_/A sky130_fd_sc_hd__or2_4
XANTENNA__18969__A _19085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15129_ _15119_/X _15129_/B _15125_/X _15128_/X VGND VGND VPWR VPWR _15130_/D sky130_fd_sc_hd__or4_4
XFILLER_126_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12082__A _12081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15845__A3 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19937_ _23575_/Q VGND VGND VPWR VPWR _19937_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22576__B1 _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19868_ _19866_/Y _19862_/X _19796_/X _19867_/X VGND VGND VPWR VPWR _19868_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12810__A _22724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22003__B _21991_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16255__B1 _15905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24688__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18819_ _18819_/A VGND VGND VPWR VPWR _18819_/Y sky130_fd_sc_hd__inv_2
XFILLER_244_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19799_ _23625_/Q VGND VGND VPWR VPWR _21899_/B sky130_fd_sc_hd__inv_2
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22328__B1 _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21830_ _21815_/A _21828_/X _21830_/C VGND VGND VPWR VPWR _21830_/X sky130_fd_sc_hd__and3_4
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24617__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12816__B1 _22678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22879__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16007__B1 _11752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21761_ _21121_/X _21759_/Y _21605_/X _21760_/X VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23115__A _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _13136_/B VGND VGND VPWR VPWR _20712_/Y sky130_fd_sc_hd__inv_2
X_23500_ _23516_/CLK _20152_/X VGND VGND VPWR VPWR _23500_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24480_ _25043_/CLK _24480_/D HRESETn VGND VGND VPWR VPWR _24480_/Q sky130_fd_sc_hd__dfrtp_4
X_21692_ _21497_/A _21692_/B VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__or2_4
XANTENNA__22954__A _24572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23553_/CLK _23431_/D VGND VGND VPWR VPWR _23431_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20643_ _17400_/X _20643_/B _20628_/X VGND VGND VPWR VPWR _20643_/X sky130_fd_sc_hd__and3_4
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14977__A1_N _15258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22673__B _22673_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _12055_/A _25175_/Q VGND VGND VPWR VPWR _23362_/X sky130_fd_sc_hd__and2_4
X_20574_ _20550_/Y VGND VGND VPWR VPWR _20574_/X sky130_fd_sc_hd__buf_2
X_22313_ _16529_/A _21450_/X _21335_/X VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__o21a_4
X_25101_ _25281_/CLK _25101_/D HRESETn VGND VGND VPWR VPWR _13577_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23293_ _24647_/Q _21536_/X VGND VGND VPWR VPWR _23293_/X sky130_fd_sc_hd__or2_4
XFILLER_192_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16730__B2 _16654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25032_ _25030_/CLK _25032_/D HRESETn VGND VGND VPWR VPWR _25032_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12347__A2 _24843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22244_ _22260_/A _22244_/B VGND VGND VPWR VPWR _22244_/X sky130_fd_sc_hd__or2_4
XFILLER_192_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20409__A3 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16089__A3 _15933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22175_ _16460_/A _22172_/X _22175_/C VGND VGND VPWR VPWR _22205_/B sky130_fd_sc_hd__and3_4
XANTENNA__12423__C _12391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21126_ _15647_/Y _21126_/B VGND VGND VPWR VPWR _21126_/X sky130_fd_sc_hd__or2_4
XFILLER_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21057_ _21047_/X _21053_/X _21882_/A _21056_/X VGND VGND VPWR VPWR _21058_/C sky130_fd_sc_hd__a211o_4
XANTENNA__19432__B1 _19341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_115_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24509_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16246__B1 _16245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20008_ _21688_/B _20006_/X _20007_/X _20006_/X VGND VGND VPWR VPWR _23551_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_178_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _25488_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_246_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12830_ _12828_/X _24794_/Q _25401_/Q _12829_/Y VGND VGND VPWR VPWR _12836_/B sky130_fd_sc_hd__a2bb2o_4
X_24816_ _24856_/CLK _24816_/D HRESETn VGND VGND VPWR VPWR _23162_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15552__A2_N _15547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21752__B _21752_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _25389_/Q VGND VGND VPWR VPWR _12762_/A sky130_fd_sc_hd__inv_2
X_24747_ _24372_/CLK _24747_/D HRESETn VGND VGND VPWR VPWR _16018_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _17727_/A _21959_/B VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__or2_4
XANTENNA__17746__B1 _21704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18119__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14499_/Y _14497_/X _14479_/X _14497_/X VGND VGND VPWR VPWR _14500_/X sky130_fd_sc_hd__a2bb2o_4
X_11712_ _11712_/A _11712_/B VGND VGND VPWR VPWR _11713_/A sky130_fd_sc_hd__and2_4
XFILLER_187_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12619_/B _12689_/B VGND VGND VPWR VPWR _12693_/C sky130_fd_sc_hd__nand2_4
X_15480_ _14400_/A VGND VGND VPWR VPWR _15480_/X sky130_fd_sc_hd__buf_2
XFILLER_188_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _24674_/CLK _16211_/X HRESETn VGND VGND VPWR VPWR _23183_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_199_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22864__A _22854_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14430_/Y _14428_/X _14400_/X _14428_/X VGND VGND VPWR VPWR _14431_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23631_/CLK _19785_/X VGND VGND VPWR VPWR _13467_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12167__A _14342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17127_/X _17143_/X _17149_/Y VGND VGND VPWR VPWR _17150_/X sky130_fd_sc_hd__and3_4
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _14362_/A VGND VGND VPWR VPWR _14362_/Y sky130_fd_sc_hd__inv_2
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _16100_/Y _16098_/X _11755_/X _16098_/X VGND VGND VPWR VPWR _16101_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13222_/X _13313_/B VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__or2_4
XFILLER_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _14293_/A VGND VGND VPWR VPWR _14293_/Y sky130_fd_sc_hd__inv_2
X_17081_ _17075_/C _17079_/A VGND VGND VPWR VPWR _17081_/X sky130_fd_sc_hd__or2_4
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13244_ _13243_/X _19679_/A VGND VGND VPWR VPWR _13244_/X sky130_fd_sc_hd__or2_4
X_16032_ _16030_/Y _16031_/X _15963_/X _16031_/X VGND VGND VPWR VPWR _24742_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _13199_/A _13175_/B VGND VGND VPWR VPWR _13176_/C sky130_fd_sc_hd__or2_4
X_12126_ _12125_/Y _12123_/X _11862_/X _12123_/X VGND VGND VPWR VPWR _12126_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15827__A3 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17983_ _18006_/A VGND VGND VPWR VPWR _17984_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19722_ _19722_/A VGND VGND VPWR VPWR _19722_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_74_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12057_ _16193_/A VGND VGND VPWR VPWR _13484_/C sky130_fd_sc_hd__buf_2
X_16934_ _24703_/Q _17832_/A _16164_/Y _16937_/A VGND VGND VPWR VPWR _16941_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19423__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19653_ _19652_/Y VGND VGND VPWR VPWR _19653_/X sky130_fd_sc_hd__buf_2
XANTENNA__24781__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16865_ _16864_/Y _16805_/X _16729_/X _16805_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11891__D _11890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18604_ _18604_/A VGND VGND VPWR VPWR _18604_/X sky130_fd_sc_hd__buf_2
XANTENNA__22758__B _22789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15816_ _15790_/X _15804_/X _15738_/X _24848_/Q _15802_/X VGND VGND VPWR VPWR _15816_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24710__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19584_ _23696_/Q VGND VGND VPWR VPWR _21828_/B sky130_fd_sc_hd__inv_2
X_16796_ _19131_/A VGND VGND VPWR VPWR _16796_/X sky130_fd_sc_hd__buf_2
XFILLER_225_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18535_ _18550_/A _18533_/X _18534_/X VGND VGND VPWR VPWR _24184_/D sky130_fd_sc_hd__and3_4
XANTENNA__24028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15747_ _12568_/Y _15744_/X _11800_/X _15744_/X VGND VGND VPWR VPWR _15747_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ _12855_/C _12958_/X _12891_/X _12955_/B VGND VGND VPWR VPWR _12959_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21533__B2 _22530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18466_ _24188_/Q VGND VGND VPWR VPWR _18467_/A sky130_fd_sc_hd__inv_2
X_15678_ _21596_/A VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__buf_2
X_17417_ _17396_/X _17410_/X _24341_/Q _21008_/A _17413_/X VGND VGND VPWR VPWR _17417_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ _14628_/Y _14629_/B _14679_/B _13547_/Y VGND VGND VPWR VPWR _14629_/X sky130_fd_sc_hd__and4_4
X_18397_ _21109_/A _17280_/X _18396_/Y VGND VGND VPWR VPWR _24195_/D sky130_fd_sc_hd__o21a_4
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17348_ _17348_/A _17348_/B VGND VGND VPWR VPWR _17350_/B sky130_fd_sc_hd__or2_4
XFILLER_228_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16922__D _16921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15388__A _15388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17279_ _17240_/X VGND VGND VPWR VPWR _17296_/A sky130_fd_sc_hd__inv_2
XANTENNA__23101__C _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12805__A _22139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19018_ _19017_/Y _19013_/X _18991_/X _19013_/X VGND VGND VPWR VPWR _23896_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20290_ _23447_/Q VGND VGND VPWR VPWR _21644_/B sky130_fd_sc_hd__inv_2
XFILLER_155_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22797__B1 _17767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24869__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21556__C _21113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23980_ _23980_/CLK _23980_/D HRESETn VGND VGND VPWR VPWR _23980_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16228__B1 _15967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22931_ _22694_/B VGND VGND VPWR VPWR _23177_/B sky130_fd_sc_hd__buf_2
XFILLER_228_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15851__A _19761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22862_ _21430_/X VGND VGND VPWR VPWR _22862_/X sky130_fd_sc_hd__buf_2
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15451__A1 _14289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24601_ _24601_/CLK _16424_/X HRESETn VGND VGND VPWR VPWR _24601_/Q sky130_fd_sc_hd__dfrtp_4
X_21813_ _21474_/A _19976_/Y VGND VGND VPWR VPWR _21815_/B sky130_fd_sc_hd__or2_4
X_22793_ _15553_/X VGND VGND VPWR VPWR _22793_/X sky130_fd_sc_hd__buf_2
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21744_ _21578_/X _21742_/X _21584_/X _21743_/X VGND VGND VPWR VPWR _21744_/X sky130_fd_sc_hd__o22a_4
X_24532_ _24532_/CLK _24532_/D HRESETn VGND VGND VPWR VPWR _16601_/A sky130_fd_sc_hd__dfrtp_4
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22684__A _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17778__A _23332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21675_/A _21675_/B VGND VGND VPWR VPWR _21677_/B sky130_fd_sc_hd__or2_4
X_24463_ _24430_/CLK _24463_/D HRESETn VGND VGND VPWR VPWR _16776_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16951__B2 _16950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20626_ _20626_/A VGND VGND VPWR VPWR _20626_/Y sky130_fd_sc_hd__inv_2
X_23414_ _23590_/CLK _20378_/X VGND VGND VPWR VPWR _23414_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24394_ _24406_/CLK _24394_/D HRESETn VGND VGND VPWR VPWR _24394_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23345_ _24616_/Q _23313_/B VGND VGND VPWR VPWR _23345_/X sky130_fd_sc_hd__or2_4
X_20557_ _18877_/X _20557_/B _20556_/X VGND VGND VPWR VPWR _20557_/X sky130_fd_sc_hd__and3_4
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23276_ _14939_/A _21551_/X _22108_/X _23275_/X VGND VGND VPWR VPWR _23277_/C sky130_fd_sc_hd__a211o_4
X_20488_ _14286_/Y _20503_/B _14290_/A VGND VGND VPWR VPWR _20535_/A sky130_fd_sc_hd__and3_4
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22227_ _22227_/A _20131_/Y VGND VGND VPWR VPWR _22228_/C sky130_fd_sc_hd__or2_4
X_25015_ _25011_/CLK _15291_/X HRESETn VGND VGND VPWR VPWR _25015_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22158_ _24726_/Q _22153_/X _22533_/A _22157_/X VGND VGND VPWR VPWR _22158_/X sky130_fd_sc_hd__a211o_4
XFILLER_160_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21109_ _21109_/A _21109_/B VGND VGND VPWR VPWR _21109_/X sky130_fd_sc_hd__and2_4
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _14980_/A VGND VGND VPWR VPWR _14980_/Y sky130_fd_sc_hd__inv_2
X_22089_ _22385_/A _20155_/Y VGND VGND VPWR VPWR _22091_/B sky130_fd_sc_hd__or2_4
XFILLER_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13931_ _13951_/A _13951_/B _13964_/A VGND VGND VPWR VPWR _13931_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_75_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15761__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _15833_/X _15652_/Y HWDATA[31] _24515_/Q _16652_/A VGND VGND VPWR VPWR _24515_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_235_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13862_ _13862_/A _13867_/A VGND VGND VPWR VPWR _13862_/Y sky130_fd_sc_hd__nor2_4
XFILLER_219_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15601_ _15601_/A VGND VGND VPWR VPWR _15601_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12813_ _12803_/X _12806_/X _12809_/X _12813_/D VGND VGND VPWR VPWR _12813_/X sky130_fd_sc_hd__or4_4
X_16581_ _24540_/Q VGND VGND VPWR VPWR _16581_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13793_ _16464_/A _16464_/B _13804_/C _13793_/D VGND VGND VPWR VPWR _13793_/X sky130_fd_sc_hd__and4_4
XFILLER_216_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18320_ _17740_/A _18319_/A _24224_/Q _21463_/A VGND VGND VPWR VPWR _18320_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13281__A _13356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15532_ _11736_/C VGND VGND VPWR VPWR _15532_/Y sky130_fd_sc_hd__inv_2
X_12744_ _12737_/B VGND VGND VPWR VPWR _12745_/B sky130_fd_sc_hd__inv_2
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18251_ _18245_/X _18247_/X _16248_/A _22631_/A _18248_/X VGND VGND VPWR VPWR _18251_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15463_ _24086_/Q _15458_/X _15450_/Y _13955_/A _15461_/X VGND VGND VPWR VPWR _24969_/D
+ sky130_fd_sc_hd__a32o_4
X_12675_ _12620_/C _12674_/X VGND VGND VPWR VPWR _12676_/B sky130_fd_sc_hd__or2_4
XANTENNA__16592__A _16618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _24636_/Q _24365_/Q _16324_/Y _17263_/C VGND VGND VPWR VPWR _17202_/X sky130_fd_sc_hd__o22a_4
XFILLER_187_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _14414_/A VGND VGND VPWR VPWR _14414_/Y sky130_fd_sc_hd__inv_2
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18182_ _17979_/A _18182_/B VGND VGND VPWR VPWR _18183_/C sky130_fd_sc_hd__or2_4
XFILLER_230_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _15137_/Y _15389_/B _15390_/Y _15348_/X VGND VGND VPWR VPWR _15394_/X sky130_fd_sc_hd__a211o_4
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11767__B1 _11766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17127_/X _17131_/X _17133_/C VGND VGND VPWR VPWR _24391_/D sky130_fd_sc_hd__and3_4
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _25171_/Q _14359_/A _14349_/D VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__and3_4
XFILLER_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17064_ _17064_/A VGND VGND VPWR VPWR _17393_/B sky130_fd_sc_hd__inv_2
X_14276_ _14275_/Y _14273_/X _13806_/X _14273_/X VGND VGND VPWR VPWR _14276_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16015_ _16014_/Y _16012_/X _15950_/X _16012_/X VGND VGND VPWR VPWR _24749_/D sky130_fd_sc_hd__a2bb2o_4
X_13227_ _13164_/Y VGND VGND VPWR VPWR _13387_/A sky130_fd_sc_hd__buf_2
XANTENNA__15936__A _15683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19644__B1 _19643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13158_ _13195_/A _13158_/B VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__or2_4
XFILLER_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12109_ _12109_/A _12107_/X _12109_/C _12108_/X VGND VGND VPWR VPWR _12110_/A sky130_fd_sc_hd__or4_4
X_13089_ _12387_/X _12342_/Y _13115_/A _13115_/B VGND VGND VPWR VPWR _13089_/X sky130_fd_sc_hd__or4_4
X_17966_ _17951_/A _18981_/A VGND VGND VPWR VPWR _17967_/C sky130_fd_sc_hd__or2_4
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16917_ _24694_/Q _24271_/Q _16156_/Y _16916_/Y VGND VGND VPWR VPWR _16922_/B sky130_fd_sc_hd__o22a_4
X_19705_ _19703_/Y _19699_/X _19659_/X _19704_/X VGND VGND VPWR VPWR _23658_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17897_ _24262_/Q VGND VGND VPWR VPWR _22009_/A sky130_fd_sc_hd__inv_2
XFILLER_226_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16767__A _16737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16848_ _14909_/Y _16846_/X _11830_/X _16846_/X VGND VGND VPWR VPWR _24429_/D sky130_fd_sc_hd__a2bb2o_4
X_19636_ _19636_/A VGND VGND VPWR VPWR _19636_/X sky130_fd_sc_hd__buf_2
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_161_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23885_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_19_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_4_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_214_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16630__B1 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19567_ _19564_/Y _19565_/X _19566_/X _19565_/X VGND VGND VPWR VPWR _19567_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_18_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _23582_/CLK sky130_fd_sc_hd__clkbuf_1
X_16779_ _16782_/A VGND VGND VPWR VPWR _16779_/X sky130_fd_sc_hd__buf_2
XFILLER_240_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22703__B1 _17766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18518_ _18467_/A _18517_/X _18494_/X VGND VGND VPWR VPWR _18518_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12798__A2 _21537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19498_ _23726_/Q VGND VGND VPWR VPWR _21501_/B sky130_fd_sc_hd__inv_2
XFILLER_178_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18449_ _24185_/Q VGND VGND VPWR VPWR _18486_/B sky130_fd_sc_hd__inv_2
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21460_ _12853_/Y _21456_/X _21459_/X VGND VGND VPWR VPWR _21460_/X sky130_fd_sc_hd__o21a_4
XFILLER_239_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20411_ _20406_/A VGND VGND VPWR VPWR _20411_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17489__A2 _17484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21391_ _21408_/A _21391_/B VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__or2_4
XFILLER_147_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23130_ _22993_/X _23128_/X _23062_/X _25550_/Q _23129_/X VGND VGND VPWR VPWR _23130_/X
+ sky130_fd_sc_hd__a32o_4
X_20342_ _20408_/A VGND VGND VPWR VPWR _20342_/X sky130_fd_sc_hd__buf_2
XFILLER_161_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23061_ _23061_/A _22882_/X VGND VGND VPWR VPWR _23061_/X sky130_fd_sc_hd__or2_4
X_20273_ _20272_/Y _20270_/X _19832_/X _20270_/X VGND VGND VPWR VPWR _23454_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12183__B1 _11871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _13826_/X VGND VGND VPWR VPWR _22595_/B sky130_fd_sc_hd__buf_2
XANTENNA__16449__B1 _16368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24632__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23963_ _23946_/CLK scl_i_S4 HRESETn VGND VGND VPWR VPWR _23964_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_229_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22942__B1 _22816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22914_ _22488_/X _22913_/X _21434_/X _24879_/Q _22784_/X VGND VGND VPWR VPWR _22914_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_217_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23894_ _24101_/CLK _19023_/X VGND VGND VPWR VPWR _19022_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_244_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16621__B1 _16537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22845_ _21295_/A VGND VGND VPWR VPWR _22845_/X sky130_fd_sc_hd__buf_2
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _22743_/X _22750_/Y _22754_/X _22775_/Y VGND VGND VPWR VPWR HRDATA[15] sky130_fd_sc_hd__or4_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20927__A _20836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24515_ _24029_/CLK _24515_/D HRESETn VGND VGND VPWR VPWR _24515_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21727_ _25110_/Q _22129_/B VGND VGND VPWR VPWR _21730_/B sky130_fd_sc_hd__nand2_4
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25495_ _24171_/CLK _25495_/D HRESETn VGND VGND VPWR VPWR _25495_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17301__A _17266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12460_ _12459_/X VGND VGND VPWR VPWR _25454_/D sky130_fd_sc_hd__inv_2
X_21658_ _21654_/X _21657_/X _25278_/Q _18268_/X VGND VGND VPWR VPWR _21658_/X sky130_fd_sc_hd__o22a_4
X_24446_ _25043_/CLK _16814_/X HRESETn VGND VGND VPWR VPWR _14914_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_184_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12391_ _12391_/A _12391_/B VGND VGND VPWR VPWR _12391_/X sky130_fd_sc_hd__or2_4
X_20609_ _20609_/A _20609_/B VGND VGND VPWR VPWR _20609_/X sky130_fd_sc_hd__or2_4
X_21589_ _15019_/Y _21589_/B VGND VGND VPWR VPWR _21589_/X sky130_fd_sc_hd__and2_4
X_24377_ _24641_/CLK _24377_/D HRESETn VGND VGND VPWR VPWR _24377_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14130_ _14414_/A _14119_/X _14120_/X _14129_/Y VGND VGND VPWR VPWR _14130_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16688__B1 _16419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23328_ _24717_/Q _23296_/B VGND VGND VPWR VPWR _23328_/X sky130_fd_sc_hd__or2_4
XFILLER_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14061_ _14024_/X _14060_/X VGND VGND VPWR VPWR _14069_/A sky130_fd_sc_hd__or2_4
XANTENNA__15756__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23259_ _23240_/X _23243_/X _23247_/Y _23258_/X VGND VGND VPWR VPWR HRDATA[28] sky130_fd_sc_hd__a211o_4
XANTENNA__14660__A _18013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13012_ _13011_/X VGND VGND VPWR VPWR _13013_/B sky130_fd_sc_hd__inv_2
XFILLER_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_6_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ _17769_/D _17820_/B VGND VGND VPWR VPWR _17820_/X sky130_fd_sc_hd__or2_4
XFILLER_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13276__A _13217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17971__A _17973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22589__A _16434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16860__B1 _16796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17751_ _17751_/A VGND VGND VPWR VPWR _17771_/A sky130_fd_sc_hd__inv_2
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14963_ _15251_/A _16841_/A _15251_/A _16841_/A VGND VGND VPWR VPWR _14972_/A sky130_fd_sc_hd__a2bb2o_4
X_16702_ _22616_/A _16697_/X _15761_/X _16697_/X VGND VGND VPWR VPWR _24495_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13914_ _13954_/B _13911_/Y _13955_/A _13913_/Y VGND VGND VPWR VPWR _13978_/B sky130_fd_sc_hd__and4_4
X_17682_ _17585_/D _17678_/X VGND VGND VPWR VPWR _17682_/Y sky130_fd_sc_hd__nand2_4
X_14894_ _25024_/Q VGND VGND VPWR VPWR _15070_/A sky130_fd_sc_hd__inv_2
XFILLER_247_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19421_ _19151_/A VGND VGND VPWR VPWR _19421_/X sky130_fd_sc_hd__buf_2
XFILLER_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16633_ _14769_/X _16184_/B _13599_/B VGND VGND VPWR VPWR _16633_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_234_0_HCLK clkbuf_8_234_0_HCLK/A VGND VGND VPWR VPWR _24095_/CLK sky130_fd_sc_hd__clkbuf_1
X_13845_ _13566_/Y _13842_/X _13844_/X _13842_/X VGND VGND VPWR VPWR _25267_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19352_ _18055_/B VGND VGND VPWR VPWR _19352_/Y sky130_fd_sc_hd__inv_2
X_16564_ _16564_/A VGND VGND VPWR VPWR _16564_/Y sky130_fd_sc_hd__inv_2
X_13776_ _13774_/X _13775_/X _13774_/X _13775_/X VGND VGND VPWR VPWR _25283_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18303_ _18297_/X _18302_/Y VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__or2_4
X_15515_ _15515_/A VGND VGND VPWR VPWR _15515_/Y sky130_fd_sc_hd__inv_2
X_12727_ _12550_/Y _12731_/A VGND VGND VPWR VPWR _12727_/Y sky130_fd_sc_hd__nand2_4
X_19283_ _19283_/A VGND VGND VPWR VPWR _19283_/Y sky130_fd_sc_hd__inv_2
X_16495_ _16495_/A VGND VGND VPWR VPWR _16495_/X sky130_fd_sc_hd__buf_2
XFILLER_231_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18234_ _18234_/A _18234_/B _18234_/C VGND VGND VPWR VPWR _18235_/C sky130_fd_sc_hd__or3_4
X_15446_ _15446_/A VGND VGND VPWR VPWR _15446_/X sky130_fd_sc_hd__buf_2
X_12658_ _12658_/A VGND VGND VPWR VPWR _25432_/D sky130_fd_sc_hd__inv_2
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18165_ _18165_/A _19180_/A VGND VGND VPWR VPWR _18166_/C sky130_fd_sc_hd__or2_4
X_15377_ _15384_/A _15377_/B _15376_/Y VGND VGND VPWR VPWR _24999_/D sky130_fd_sc_hd__and3_4
XFILLER_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12589_ _12588_/Y _12595_/A _12622_/A _12532_/Y VGND VGND VPWR VPWR _12589_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _16996_/Y _17119_/B VGND VGND VPWR VPWR _17117_/C sky130_fd_sc_hd__nand2_4
X_14328_ _25178_/Q _14308_/Y _25177_/Q _14316_/A VGND VGND VPWR VPWR _14328_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21668__A _21668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18096_ _18131_/A _18096_/B _18095_/X VGND VGND VPWR VPWR _18107_/B sky130_fd_sc_hd__or3_4
XFILLER_128_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17047_ _16992_/Y _17142_/A _16987_/Y _16969_/Y VGND VGND VPWR VPWR _17047_/X sky130_fd_sc_hd__or4_4
X_14259_ _14259_/A _13953_/Y _13968_/Y VGND VGND VPWR VPWR _14260_/D sky130_fd_sc_hd__or3_4
XANTENNA__18042__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12165__B1 _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20227__B2 _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18998_ _23901_/Q VGND VGND VPWR VPWR _18998_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16851__B1 _16613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_44_0_HCLK clkbuf_6_44_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17945_/A _17947_/X _17948_/X VGND VGND VPWR VPWR _17949_/X sky130_fd_sc_hd__and3_4
XFILLER_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16497__A _24572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20960_ _13676_/A VGND VGND VPWR VPWR _20960_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15406__A1 _15082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19619_ _23685_/Q VGND VGND VPWR VPWR _19619_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20891_ _13672_/A VGND VGND VPWR VPWR _20891_/Y sky130_fd_sc_hd__inv_2
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22630_ _13555_/Y _22706_/B VGND VGND VPWR VPWR _22630_/X sky130_fd_sc_hd__and2_4
XFILLER_41_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22152__A1 _24351_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ _22754_/A _22561_/B _22561_/C VGND VGND VPWR VPWR _22588_/C sky130_fd_sc_hd__and3_4
XANTENNA__23123__A _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21512_ _21487_/X _21509_/X _21511_/X VGND VGND VPWR VPWR _21512_/Y sky130_fd_sc_hd__a21oi_4
X_24300_ _24937_/CLK _24300_/D HRESETn VGND VGND VPWR VPWR _24300_/Q sky130_fd_sc_hd__dfrtp_4
X_22492_ _22430_/A _22492_/B VGND VGND VPWR VPWR _22506_/C sky130_fd_sc_hd__and2_4
X_25280_ _23647_/CLK _13807_/X HRESETn VGND VGND VPWR VPWR _13795_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21443_ _21543_/A VGND VGND VPWR VPWR _23016_/A sky130_fd_sc_hd__buf_2
X_24231_ _24238_/CLK _24231_/D HRESETn VGND VGND VPWR VPWR _24231_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24162_ _25212_/CLK _18709_/X HRESETn VGND VGND VPWR VPWR _24162_/Q sky130_fd_sc_hd__dfrtp_4
X_21374_ _21372_/Y _21161_/X _17443_/Y _21733_/B VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24884__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20325_ _22365_/B _20324_/X _19990_/X _20324_/X VGND VGND VPWR VPWR _23435_/D sky130_fd_sc_hd__a2bb2o_4
X_23113_ _21126_/B VGND VGND VPWR VPWR _23113_/X sky130_fd_sc_hd__buf_2
XFILLER_134_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24093_ _23980_/CLK _20512_/X HRESETn VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19048__A _19048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24813__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23044_ _16120_/Y _22531_/B _22861_/X _11782_/Y _22864_/X VGND VGND VPWR VPWR _23044_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_190_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_126_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20256_ _24213_/Q _18342_/A _20079_/A _20256_/D VGND VGND VPWR VPWR _20256_/X sky130_fd_sc_hd__or4_4
XFILLER_150_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20187_ _21407_/B _20184_/X _20122_/X _20184_/X VGND VGND VPWR VPWR _20187_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16842__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24995_ _24981_/CLK _15386_/Y HRESETn VGND VGND VPWR VPWR _15139_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22202__A _21877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11960_ _19646_/A VGND VGND VPWR VPWR _11960_/Y sky130_fd_sc_hd__inv_2
X_23946_ _23946_/CLK _20993_/X HRESETn VGND VGND VPWR VPWR _20994_/A sky130_fd_sc_hd__dfstp_4
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11891_ _25524_/Q _11897_/A _11879_/A _11890_/X VGND VGND VPWR VPWR _11891_/X sky130_fd_sc_hd__and4_4
X_23877_ _24214_/CLK _23877_/D VGND VGND VPWR VPWR _19072_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_244_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13630_ _13628_/A _13628_/B _14670_/A VGND VGND VPWR VPWR _13630_/X sky130_fd_sc_hd__a21o_4
XFILLER_204_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22828_ _22854_/B VGND VGND VPWR VPWR _22954_/B sky130_fd_sc_hd__buf_2
XFILLER_204_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_64_0_HCLK clkbuf_7_32_0_HCLK/X VGND VGND VPWR VPWR _24283_/CLK sky130_fd_sc_hd__clkbuf_1
X_13561_ _13561_/A VGND VGND VPWR VPWR _13561_/Y sky130_fd_sc_hd__inv_2
X_25547_ _24327_/CLK _25547_/D HRESETn VGND VGND VPWR VPWR _25547_/Q sky130_fd_sc_hd__dfrtp_4
X_22759_ _22494_/X _22758_/X _21303_/A _24840_/Q _22498_/X VGND VGND VPWR VPWR _22759_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14655__A _18097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15300_ _15299_/Y VGND VGND VPWR VPWR _15388_/A sky130_fd_sc_hd__buf_2
XFILLER_158_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12512_ _12501_/A _12508_/X _12512_/C VGND VGND VPWR VPWR _25440_/D sky130_fd_sc_hd__and3_4
X_16280_ _16280_/A _16001_/X VGND VGND VPWR VPWR _16280_/X sky130_fd_sc_hd__or2_4
X_13492_ _13490_/Y _13486_/X _11851_/X _13491_/X VGND VGND VPWR VPWR _25327_/D sky130_fd_sc_hd__a2bb2o_4
X_25478_ _24119_/CLK _12124_/X HRESETn VGND VGND VPWR VPWR _12122_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22872__A _22157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15231_ _15231_/A _15219_/X VGND VGND VPWR VPWR _15231_/X sky130_fd_sc_hd__or2_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _12442_/X VGND VGND VPWR VPWR _12444_/B sky130_fd_sc_hd__inv_2
X_24429_ _24430_/CLK _24429_/D HRESETn VGND VGND VPWR VPWR _14909_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12175__A _12175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15162_ _15162_/A VGND VGND VPWR VPWR _15162_/Y sky130_fd_sc_hd__inv_2
X_12374_ _13004_/B _24829_/Q _12994_/A _12373_/Y VGND VGND VPWR VPWR _12374_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14113_ _14112_/X VGND VGND VPWR VPWR _14115_/B sky130_fd_sc_hd__inv_2
XFILLER_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24554__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15093_ _15092_/Y VGND VGND VPWR VPWR _15380_/A sky130_fd_sc_hd__buf_2
X_19970_ _19969_/Y _19967_/X _19629_/X _19967_/X VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14390__A _14116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14044_ _14043_/X VGND VGND VPWR VPWR _14045_/C sky130_fd_sc_hd__inv_2
X_18921_ _23930_/Q VGND VGND VPWR VPWR _22080_/B sky130_fd_sc_hd__inv_2
XFILLER_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18852_ _24557_/Q _18809_/A _16522_/A _18794_/C VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17803_ _17771_/A _17802_/X VGND VGND VPWR VPWR _17803_/X sky130_fd_sc_hd__or2_4
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18783_ _18699_/A _18780_/X VGND VGND VPWR VPWR _18784_/C sky130_fd_sc_hd__or2_4
X_15995_ _15486_/A VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__buf_2
XFILLER_95_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17734_ _17733_/X VGND VGND VPWR VPWR _17734_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14946_ _24421_/Q VGND VGND VPWR VPWR _14946_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21951__A _21679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17665_ _17667_/B VGND VGND VPWR VPWR _17666_/B sky130_fd_sc_hd__inv_2
XFILLER_236_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14877_ _24958_/Q VGND VGND VPWR VPWR _14877_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16616_ _16615_/Y _16610_/X _16530_/X _16610_/X VGND VGND VPWR VPWR _16616_/X sky130_fd_sc_hd__a2bb2o_4
X_19404_ _18143_/B VGND VGND VPWR VPWR _19404_/Y sky130_fd_sc_hd__inv_2
X_13828_ _13781_/A _13782_/A _13828_/C _13828_/D VGND VGND VPWR VPWR _13828_/X sky130_fd_sc_hd__and4_4
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19421__A _19151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17596_ _17596_/A _17596_/B VGND VGND VPWR VPWR _17598_/B sky130_fd_sc_hd__or2_4
XFILLER_223_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16547_ _16546_/Y _16469_/X _16276_/X _16469_/X VGND VGND VPWR VPWR _24553_/D sky130_fd_sc_hd__a2bb2o_4
X_19335_ _23784_/Q VGND VGND VPWR VPWR _19335_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13759_ _25282_/Q VGND VGND VPWR VPWR _13759_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22685__A2 _23027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19266_ _23809_/Q VGND VGND VPWR VPWR _21896_/B sky130_fd_sc_hd__inv_2
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16478_ _16478_/A VGND VGND VPWR VPWR _16478_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18217_ _18084_/X _23901_/Q VGND VGND VPWR VPWR _18217_/X sky130_fd_sc_hd__or2_4
X_15429_ _15424_/X _15429_/B _15427_/C VGND VGND VPWR VPWR _15429_/X sky130_fd_sc_hd__and3_4
X_19197_ _19195_/Y _19191_/X _19151_/X _19196_/X VGND VGND VPWR VPWR _19197_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18148_ _18051_/A _18144_/X _18148_/C VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__or3_4
XFILLER_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18079_ _18227_/A _18075_/X _18078_/X VGND VGND VPWR VPWR _18079_/X sky130_fd_sc_hd__or3_4
X_20110_ _20107_/Y _20101_/X _20108_/X _20109_/X VGND VGND VPWR VPWR _20110_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _21090_/A VGND VGND VPWR VPWR _21091_/B sky130_fd_sc_hd__buf_2
X_20041_ _23539_/Q VGND VGND VPWR VPWR _22271_/B sky130_fd_sc_hd__inv_2
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17550__A1_N _11853_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16824__B1 HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23118__A _21535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23800_ _23529_/CLK _23800_/D VGND VGND VPWR VPWR _23800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24780_ _24781_/CLK _15954_/X HRESETn VGND VGND VPWR VPWR _23196_/A sky130_fd_sc_hd__dfrtp_4
X_21992_ _18366_/Y _23423_/Q _24206_/Q _20356_/Y VGND VGND VPWR VPWR _21992_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21176__A2 _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _23555_/CLK _19487_/X VGND VGND VPWR VPWR _23731_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _20944_/A VGND VGND VPWR VPWR _20943_/Y sky130_fd_sc_hd__inv_2
XPHY_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23654_/CLK _23662_/D VGND VGND VPWR VPWR _23662_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _24056_/Q VGND VGND VPWR VPWR _20874_/Y sky130_fd_sc_hd__inv_2
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25401_ _25402_/CLK _25401_/D HRESETn VGND VGND VPWR VPWR _25401_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _22613_/A _21103_/A VGND VGND VPWR VPWR _22613_/X sky130_fd_sc_hd__or2_4
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23593_ _23684_/CLK _23593_/D VGND VGND VPWR VPWR _19890_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__14475__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13810__B1 _13809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20687__A1 _20681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25332_ _25488_/CLK _25332_/D HRESETn VGND VGND VPWR VPWR _25332_/Q sky130_fd_sc_hd__dfrtp_4
X_22544_ _23148_/A VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__buf_2
XFILLER_194_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25263_ _25276_/CLK _13853_/X HRESETn VGND VGND VPWR VPWR _25263_/Q sky130_fd_sc_hd__dfrtp_4
X_22475_ _20870_/C _23144_/A _16708_/Y _22289_/X VGND VGND VPWR VPWR _22476_/B sky130_fd_sc_hd__o22a_4
XFILLER_194_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24214_ _24214_/CLK _24214_/D HRESETn VGND VGND VPWR VPWR _18332_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21426_ _21605_/A VGND VGND VPWR VPWR _21427_/A sky130_fd_sc_hd__buf_2
X_25194_ _25253_/CLK _14276_/X HRESETn VGND VGND VPWR VPWR _25194_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21100__A2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21101__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21357_ _14437_/Y _21356_/X _14477_/Y _17424_/A VGND VGND VPWR VPWR _21357_/X sky130_fd_sc_hd__o22a_4
X_24145_ _24145_/CLK _24145_/D HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12129__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20308_ _20302_/Y VGND VGND VPWR VPWR _20308_/X sky130_fd_sc_hd__buf_2
X_12090_ _12090_/A VGND VGND VPWR VPWR _12090_/Y sky130_fd_sc_hd__inv_2
X_21288_ _22523_/A VGND VGND VPWR VPWR _21288_/X sky130_fd_sc_hd__buf_2
X_24076_ _24073_/CLK _24076_/D HRESETn VGND VGND VPWR VPWR _13676_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_150_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20239_ _23466_/Q VGND VGND VPWR VPWR _20239_/Y sky130_fd_sc_hd__inv_2
X_23027_ _16317_/A _23027_/B _22830_/C VGND VGND VPWR VPWR _23027_/X sky130_fd_sc_hd__and3_4
XANTENNA__13847__A1_N _13560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16144__A1_N _16143_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14800_ _19346_/A _14799_/X _19346_/A _14799_/X VGND VGND VPWR VPWR _14801_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23333__A1_N _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15780_ _12571_/Y _15772_/X _14479_/X _15726_/X VGND VGND VPWR VPWR _15780_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12992_ _24786_/Q VGND VGND VPWR VPWR _12992_/Y sky130_fd_sc_hd__inv_2
X_24978_ _24979_/CLK _15449_/X HRESETn VGND VGND VPWR VPWR _24978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14731_ _14717_/X _14730_/X VGND VGND VPWR VPWR _14731_/X sky130_fd_sc_hd__or2_4
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11943_ _19629_/A VGND VGND VPWR VPWR _11943_/X sky130_fd_sc_hd__buf_2
X_23929_ _23577_/CLK _18925_/X VGND VGND VPWR VPWR _23929_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20375__B1 _19639_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17450_ _14232_/B _17450_/B VGND VGND VPWR VPWR _17450_/Y sky130_fd_sc_hd__nor2_4
X_14662_ _17951_/A _14652_/Y VGND VGND VPWR VPWR _14662_/X sky130_fd_sc_hd__or2_4
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11874_ HWDATA[0] VGND VGND VPWR VPWR _13818_/A sky130_fd_sc_hd__buf_2
X_16401_ _16400_/Y _16398_/X _16309_/X _16398_/X VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22116__B2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13613_ _13613_/A _13613_/B VGND VGND VPWR VPWR _13614_/B sky130_fd_sc_hd__and2_4
X_17381_ _24351_/Q _17380_/Y VGND VGND VPWR VPWR _17381_/X sky130_fd_sc_hd__or2_4
X_14593_ _14593_/A _14582_/Y VGND VGND VPWR VPWR _14593_/X sky130_fd_sc_hd__or2_4
X_19120_ _19119_/X VGND VGND VPWR VPWR _19134_/A sky130_fd_sc_hd__inv_2
XFILLER_41_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16332_ _16290_/A VGND VGND VPWR VPWR _16352_/A sky130_fd_sc_hd__buf_2
XFILLER_201_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13544_ SSn_S2 _13543_/Y _13524_/X _13543_/Y VGND VGND VPWR VPWR _25309_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19051_ _19050_/Y _19044_/X _18999_/X _19037_/A VGND VGND VPWR VPWR _19051_/X sky130_fd_sc_hd__a2bb2o_4
X_16263_ _16263_/A VGND VGND VPWR VPWR _16263_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24735__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13475_ _11721_/A VGND VGND VPWR VPWR _16378_/B sky130_fd_sc_hd__buf_2
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_8_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18002_ _18191_/A _18002_/B _18002_/C VGND VGND VPWR VPWR _18003_/C sky130_fd_sc_hd__and3_4
X_15214_ _15078_/X _15181_/B _15009_/X VGND VGND VPWR VPWR _15215_/C sky130_fd_sc_hd__o21a_4
X_12426_ _12428_/B VGND VGND VPWR VPWR _12427_/B sky130_fd_sc_hd__inv_2
X_16194_ _16193_/X VGND VGND VPWR VPWR _16468_/B sky130_fd_sc_hd__buf_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23092__A2 _21039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19296__B2 _19293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15145_ _15346_/A _24608_/Q _15346_/A _24608_/Q VGND VGND VPWR VPWR _15145_/X sky130_fd_sc_hd__a2bb2o_4
X_12357_ _13006_/B _24837_/Q _13006_/B _24837_/Q VGND VGND VPWR VPWR _12357_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15857__A1 _15678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15076_ _14921_/A _15232_/A _15076_/C _14906_/Y VGND VGND VPWR VPWR _15077_/D sky130_fd_sc_hd__or4_4
X_19953_ _19953_/A VGND VGND VPWR VPWR _19953_/Y sky130_fd_sc_hd__inv_2
X_12288_ _25448_/Q VGND VGND VPWR VPWR _12288_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14027_ _14027_/A _14027_/B _14027_/C _14027_/D VGND VGND VPWR VPWR _14545_/A sky130_fd_sc_hd__or4_4
X_18904_ _23934_/Q VGND VGND VPWR VPWR _18904_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19884_ _22346_/B _19883_/X _19626_/X _19883_/X VGND VGND VPWR VPWR _23596_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18835_ _18831_/X _18832_/X _18833_/X _18834_/X VGND VGND VPWR VPWR _18851_/A sky130_fd_sc_hd__or4_4
XFILLER_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15978_ _15974_/X _15977_/X _16238_/A _22758_/A _15975_/X VGND VGND VPWR VPWR _24768_/D
+ sky130_fd_sc_hd__a32o_4
X_18766_ _18776_/A _18766_/B _18765_/Y VGND VGND VPWR VPWR _24149_/D sky130_fd_sc_hd__and3_4
XANTENNA__22777__A _21126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14929_ _14927_/A _24443_/Q _15203_/A _14928_/Y VGND VGND VPWR VPWR _14929_/X sky130_fd_sc_hd__o22a_4
X_17717_ _24222_/Q VGND VGND VPWR VPWR _17717_/X sky130_fd_sc_hd__buf_2
XFILLER_36_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18697_ _24147_/Q VGND VGND VPWR VPWR _18763_/A sky130_fd_sc_hd__inv_2
XFILLER_222_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12843__B2 _21712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22496__B _22789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19151__A _19151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17648_ _17516_/Y _17652_/B _17647_/Y VGND VGND VPWR VPWR _17648_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17579_ _17579_/A _17579_/B _17579_/C VGND VGND VPWR VPWR _17621_/D sky130_fd_sc_hd__or3_4
XANTENNA__22658__A2 _22678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19318_ _13428_/B VGND VGND VPWR VPWR _19318_/Y sky130_fd_sc_hd__inv_2
X_20590_ _14434_/Y _20574_/X _20564_/X _20589_/X VGND VGND VPWR VPWR _20591_/A sky130_fd_sc_hd__a211o_4
XFILLER_32_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _19249_/A VGND VGND VPWR VPWR _19249_/X sky130_fd_sc_hd__buf_2
XFILLER_149_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15545__B1 HADDR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22260_ _22260_/A _20367_/Y VGND VGND VPWR VPWR _22262_/B sky130_fd_sc_hd__or2_4
XFILLER_164_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19287__B2 _19286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21211_ _21211_/A _21211_/B VGND VGND VPWR VPWR _21212_/C sky130_fd_sc_hd__or2_4
XFILLER_145_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22191_ _15474_/Y _21370_/X _14235_/Y _21356_/X VGND VGND VPWR VPWR _22192_/A sky130_fd_sc_hd__o22a_4
XFILLER_133_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18495__C1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21142_ _14501_/Y _21375_/A _14191_/Y _14443_/A VGND VGND VPWR VPWR _21143_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18863__A1_N _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21073_ _21073_/A VGND VGND VPWR VPWR _21073_/Y sky130_fd_sc_hd__inv_2
X_20024_ _20024_/A VGND VGND VPWR VPWR _21944_/B sky130_fd_sc_hd__inv_2
X_24901_ _24485_/CLK _15642_/X HRESETn VGND VGND VPWR VPWR _24901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24832_ _24849_/CLK _24832_/D HRESETn VGND VGND VPWR VPWR _24832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_227_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24763_ _24759_/CLK _24763_/D HRESETn VGND VGND VPWR VPWR _22568_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20357__B1 _20249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _14626_/A _19619_/Y _14624_/A _21976_/B VGND VGND VPWR VPWR _21975_/X sky130_fd_sc_hd__o22a_4
XPHY_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23714_ _23408_/CLK _19535_/X VGND VGND VPWR VPWR _19533_/A sky130_fd_sc_hd__dfxtp_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _20900_/X _20925_/Y _24504_/Q _20904_/X VGND VGND VPWR VPWR _24067_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24694_ _25444_/CLK _24694_/D HRESETn VGND VGND VPWR VPWR _24694_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18970__B1 _18969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23647_/CLK _23645_/D VGND VGND VPWR VPWR _13464_/B sky130_fd_sc_hd__dfxtp_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12840__A2_N _23290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _16715_/Y _20854_/X _20842_/X _20856_/X VGND VGND VPWR VPWR _20858_/A sky130_fd_sc_hd__o22a_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23576_ _23488_/CLK _19936_/X VGND VGND VPWR VPWR _23576_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _20788_/A VGND VGND VPWR VPWR _20788_/X sky130_fd_sc_hd__buf_2
XANTENNA__18722__B1 _18714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25315_ _25188_/CLK _25315_/D HRESETn VGND VGND VPWR VPWR _25315_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22527_ _22527_/A _13792_/A _21383_/A VGND VGND VPWR VPWR _22527_/X sky130_fd_sc_hd__or3_4
XANTENNA__15536__B1 HADDR[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_138_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _25077_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13260_ _13178_/A _13260_/B VGND VGND VPWR VPWR _13260_/X sky130_fd_sc_hd__or2_4
X_25246_ _25246_/CLK _14076_/X HRESETn VGND VGND VPWR VPWR _25246_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22458_ _22454_/X _22458_/B _22510_/C VGND VGND VPWR VPWR _22458_/X sky130_fd_sc_hd__or3_4
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15152__A2_N _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ _25446_/Q VGND VGND VPWR VPWR _12212_/A sky130_fd_sc_hd__inv_2
XANTENNA__17289__B1 _17288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21409_ _14700_/X _21407_/X _21409_/C VGND VGND VPWR VPWR _21409_/X sky130_fd_sc_hd__and3_4
X_13191_ _13195_/A _19232_/A VGND VGND VPWR VPWR _13193_/B sky130_fd_sc_hd__or2_4
X_25177_ _25177_/CLK _14331_/X HRESETn VGND VGND VPWR VPWR _25177_/Q sky130_fd_sc_hd__dfrtp_4
X_22389_ _22090_/A _20099_/Y VGND VGND VPWR VPWR _22390_/C sky130_fd_sc_hd__or2_4
XANTENNA__22821__A2 _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12142_ _24113_/Q _12134_/B _12141_/Y VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__o21a_4
X_24128_ _23946_/CLK _18895_/X HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17963__B _17963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12073_ _12073_/A VGND VGND VPWR VPWR _13821_/B sky130_fd_sc_hd__buf_2
X_16950_ _16950_/A VGND VGND VPWR VPWR _16950_/Y sky130_fd_sc_hd__inv_2
X_24059_ _24532_/CLK _20890_/X HRESETn VGND VGND VPWR VPWR _13671_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22585__A1 _12855_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15901_ _15894_/X _15895_/X _16248_/A _22641_/A _15896_/X VGND VGND VPWR VPWR _15901_/X
+ sky130_fd_sc_hd__a32o_4
X_16881_ _16874_/X VGND VGND VPWR VPWR _16881_/X sky130_fd_sc_hd__buf_2
XFILLER_238_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15832_ _15825_/X _15828_/X _15759_/X _24837_/Q _15826_/X VGND VGND VPWR VPWR _15832_/X
+ sky130_fd_sc_hd__a32o_4
X_18620_ _16578_/A _18756_/A _16564_/A _18703_/A VGND VGND VPWR VPWR _18623_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15763_ _15772_/A VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__buf_2
X_18551_ _18539_/B VGND VGND VPWR VPWR _18552_/B sky130_fd_sc_hd__inv_2
X_12975_ _25378_/Q _12974_/Y VGND VGND VPWR VPWR _12975_/X sky130_fd_sc_hd__or2_4
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14714_ _13753_/X _14713_/Y VGND VGND VPWR VPWR _14714_/X sky130_fd_sc_hd__or2_4
X_17502_ _11824_/Y _24307_/Q _11824_/Y _24307_/Q VGND VGND VPWR VPWR _17507_/A sky130_fd_sc_hd__a2bb2o_4
X_11926_ _11885_/X _11910_/X VGND VGND VPWR VPWR _11926_/Y sky130_fd_sc_hd__nor2_4
X_18482_ _18482_/A _18480_/Y _18433_/Y _18565_/B VGND VGND VPWR VPWR _18482_/X sky130_fd_sc_hd__or4_4
X_15694_ _15701_/B VGND VGND VPWR VPWR _15694_/X sky130_fd_sc_hd__buf_2
XANTENNA__24987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17433_ _14427_/A VGND VGND VPWR VPWR _17433_/X sky130_fd_sc_hd__buf_2
XFILLER_178_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14645_ _18089_/A VGND VGND VPWR VPWR _18069_/A sky130_fd_sc_hd__buf_2
XANTENNA__21006__A scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11857_ _11749_/X VGND VGND VPWR VPWR _11857_/X sky130_fd_sc_hd__buf_2
XANTENNA__24916__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ _17364_/A _17364_/B _17364_/C VGND VGND VPWR VPWR _17364_/X sky130_fd_sc_hd__or3_4
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14576_ _14603_/A _14575_/X VGND VGND VPWR VPWR _14577_/B sky130_fd_sc_hd__or2_4
XANTENNA__23210__A1_N _17294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ _11785_/Y _11786_/X _11787_/X _11786_/X VGND VGND VPWR VPWR _25546_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_34_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_34_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16315_ HWDATA[23] VGND VGND VPWR VPWR _16315_/X sky130_fd_sc_hd__buf_2
X_19103_ _19102_/Y _19100_/X _16876_/X _19100_/X VGND VGND VPWR VPWR _23867_/D sky130_fd_sc_hd__a2bb2o_4
X_13527_ _13526_/Y _13521_/X _13481_/X _13521_/X VGND VGND VPWR VPWR _25312_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15939__A _15793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15527__B1 HADDR[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_97_0_HCLK clkbuf_7_97_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17295_ _17242_/X _17295_/B _17295_/C VGND VGND VPWR VPWR _24373_/D sky130_fd_sc_hd__and3_4
XFILLER_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19034_ _19034_/A VGND VGND VPWR VPWR _19034_/Y sky130_fd_sc_hd__inv_2
X_16246_ _16244_/Y _16242_/X _16245_/X _16242_/X VGND VGND VPWR VPWR _16246_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13458_ _13282_/A _13458_/B VGND VGND VPWR VPWR _13458_/X sky130_fd_sc_hd__or2_4
XANTENNA__14562__B HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12409_ _12225_/Y _12409_/B VGND VGND VPWR VPWR _12409_/X sky130_fd_sc_hd__or2_4
XANTENNA__13459__A _13322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16177_ _14789_/Y _14773_/Y VGND VGND VPWR VPWR _16185_/A sky130_fd_sc_hd__and2_4
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13389_ _13421_/A _23519_/Q VGND VGND VPWR VPWR _13390_/C sky130_fd_sc_hd__or2_4
XFILLER_115_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15128_ _24999_/Q _24603_/Q _15376_/A _15127_/Y VGND VGND VPWR VPWR _15128_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21676__A _21676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15674__A _15674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15059_ _14910_/Y _24477_/Q _15075_/D _24471_/Q VGND VGND VPWR VPWR _15059_/X sky130_fd_sc_hd__a2bb2o_4
X_19936_ _21780_/B _19931_/X _19803_/X _19931_/X VGND VGND VPWR VPWR _19936_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14502__B2 _14485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22576__B2 _22940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19867_ _19861_/Y VGND VGND VPWR VPWR _19867_/X sky130_fd_sc_hd__buf_2
XFILLER_110_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18818_ _18685_/Y _18791_/X _18729_/X _18815_/Y VGND VGND VPWR VPWR _18819_/A sky130_fd_sc_hd__a211o_4
X_19798_ _22072_/B _19789_/X _19796_/X _19797_/X VGND VGND VPWR VPWR _23626_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_244_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22328__B2 _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18749_ _18749_/A VGND VGND VPWR VPWR _18776_/A sky130_fd_sc_hd__buf_2
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21760_ _20846_/Y _21606_/X _24018_/Q _21607_/X VGND VGND VPWR VPWR _21760_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20711_ _20711_/A VGND VGND VPWR VPWR _20711_/Y sky130_fd_sc_hd__inv_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15766__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24657__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21691_ _21466_/X _21691_/B VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__or2_4
XANTENNA__22954__B _22954_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23430_ _23534_/CLK _23430_/D VGND VGND VPWR VPWR _20335_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20642_ _17400_/A _17399_/X VGND VGND VPWR VPWR _20643_/B sky130_fd_sc_hd__nand2_4
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20573_ _20573_/A VGND VGND VPWR VPWR _23953_/D sky130_fd_sc_hd__inv_2
X_23361_ _13474_/A _25302_/Q VGND VGND VPWR VPWR _23361_/X sky130_fd_sc_hd__and2_4
XFILLER_149_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15518__B1 HADDR[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25100_ _25281_/CLK _25100_/D HRESETn VGND VGND VPWR VPWR _14567_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22312_ _22312_/A _22945_/A VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__or2_4
XFILLER_192_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23292_ _23118_/X _23292_/B VGND VGND VPWR VPWR _23299_/C sky130_fd_sc_hd__and2_4
XFILLER_164_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22970__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20144__A2_N _20141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25031_ _25030_/CLK _15234_/X HRESETn VGND VGND VPWR VPWR _14920_/A sky130_fd_sc_hd__dfrtp_4
X_22243_ _21210_/A VGND VGND VPWR VPWR _22260_/A sky130_fd_sc_hd__buf_2
XFILLER_180_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12752__B1 _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22174_ _16617_/A _21341_/X _15676_/A _22173_/X VGND VGND VPWR VPWR _22175_/C sky130_fd_sc_hd__a211o_4
XFILLER_132_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15584__A _15584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21125_ _21231_/A VGND VGND VPWR VPWR _21126_/B sky130_fd_sc_hd__buf_2
XFILLER_160_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20159__A2_N _20156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21056_ _21056_/A _21109_/B VGND VGND VPWR VPWR _21056_/X sky130_fd_sc_hd__and2_4
XFILLER_101_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20007_ _20007_/A VGND VGND VPWR VPWR _20007_/X sky130_fd_sc_hd__buf_2
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24815_ _24883_/CLK _24815_/D HRESETn VGND VGND VPWR VPWR _23119_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12760_ _12752_/X _12760_/B _12760_/C _12760_/D VGND VGND VPWR VPWR _12800_/A sky130_fd_sc_hd__or4_4
X_24746_ _24372_/CLK _24746_/D HRESETn VGND VGND VPWR VPWR _16021_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _21954_/X _21957_/X _17732_/A VGND VGND VPWR VPWR _21966_/B sky130_fd_sc_hd__o21a_4
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17746__A1 _17710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18943__B1 _17430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _25506_/Q _25505_/Q _25507_/Q VGND VGND VPWR VPWR _11712_/B sky130_fd_sc_hd__and3_4
XFILLER_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20900_/X _20908_/X _16689_/A _20904_/X VGND VGND VPWR VPWR _20909_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15757__B1 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12680_/A _12691_/B _12690_/Y VGND VGND VPWR VPWR _25424_/D sky130_fd_sc_hd__and3_4
X_24677_ _24674_/CLK _16213_/X HRESETn VGND VGND VPWR VPWR _16212_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _22430_/A _21883_/X _21101_/X _21888_/X VGND VGND VPWR VPWR _21893_/A sky130_fd_sc_hd__a211o_4
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A VGND VGND VPWR VPWR _14430_/Y sky130_fd_sc_hd__inv_2
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _23628_/CLK _23628_/D VGND VGND VPWR VPWR _23628_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_202_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _14349_/C _14349_/D _14334_/X _14360_/X VGND VGND VPWR VPWR _14362_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15759__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15509__B1 HADDR[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23559_ _24937_/CLK _23559_/D VGND VGND VPWR VPWR _19978_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_52_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _23296_/A VGND VGND VPWR VPWR _16100_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13413_/A _13312_/B VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__or2_4
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _17080_/A _17080_/B VGND VGND VPWR VPWR _17082_/B sky130_fd_sc_hd__or2_4
XFILLER_167_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14292_ _13893_/X _20684_/A _13893_/X _14291_/X VGND VGND VPWR VPWR _14293_/A sky130_fd_sc_hd__o22a_4
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16031_ _16019_/A VGND VGND VPWR VPWR _16031_/X sky130_fd_sc_hd__buf_2
X_13243_ _13155_/X VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__buf_2
X_25229_ _23395_/CLK _14140_/X HRESETn VGND VGND VPWR VPWR _25229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21496__A _22271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13174_ _13192_/A VGND VGND VPWR VPWR _13199_/A sky130_fd_sc_hd__buf_2
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12125_ _12125_/A VGND VGND VPWR VPWR _12125_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15494__A HTRANS[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17982_ _13613_/B VGND VGND VPWR VPWR _18006_/A sky130_fd_sc_hd__buf_2
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12911__A _22678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19721_ _19717_/Y _19720_/X _19677_/X _19720_/X VGND VGND VPWR VPWR _23652_/D sky130_fd_sc_hd__a2bb2o_4
X_12056_ _14199_/A VGND VGND VPWR VPWR _16193_/A sky130_fd_sc_hd__buf_2
X_16933_ _16933_/A VGND VGND VPWR VPWR _17832_/A sky130_fd_sc_hd__inv_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19652_ _19652_/A VGND VGND VPWR VPWR _19652_/Y sky130_fd_sc_hd__inv_2
X_16864_ _24419_/Q VGND VGND VPWR VPWR _16864_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18603_ _18603_/A VGND VGND VPWR VPWR _18603_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15815_ _12330_/Y _15811_/X _11776_/X _15811_/X VGND VGND VPWR VPWR _24849_/D sky130_fd_sc_hd__a2bb2o_4
X_16795_ HWDATA[3] VGND VGND VPWR VPWR _19131_/A sky130_fd_sc_hd__buf_2
X_19583_ _21962_/B _19580_/X _11952_/X _19580_/X VGND VGND VPWR VPWR _19583_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15996__B1 _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19187__B1 _19139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15746_ _12564_/Y _15744_/X _11797_/X _15744_/X VGND VGND VPWR VPWR _15746_/X sky130_fd_sc_hd__a2bb2o_4
X_18534_ _18534_/A _18534_/B VGND VGND VPWR VPWR _18534_/X sky130_fd_sc_hd__or2_4
X_12958_ _12855_/A _12777_/X _12952_/X VGND VGND VPWR VPWR _12958_/X sky130_fd_sc_hd__or3_4
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11909_ _17711_/A _11880_/Y VGND VGND VPWR VPWR _11910_/A sky130_fd_sc_hd__and2_4
XANTENNA__24750__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15677_ _15676_/X VGND VGND VPWR VPWR _21596_/A sky130_fd_sc_hd__buf_2
X_18465_ _24186_/Q VGND VGND VPWR VPWR _18516_/A sky130_fd_sc_hd__inv_2
XFILLER_206_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12889_ _12864_/A _12886_/X VGND VGND VPWR VPWR _12889_/X sky130_fd_sc_hd__or2_4
X_14628_ _13601_/A VGND VGND VPWR VPWR _14628_/Y sky130_fd_sc_hd__inv_2
X_17416_ _17396_/X _17410_/X _24004_/Q _24343_/Q _17413_/X VGND VGND VPWR VPWR _24343_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18396_ _24649_/Q VGND VGND VPWR VPWR _18396_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17347_ _17347_/A VGND VGND VPWR VPWR _17348_/B sky130_fd_sc_hd__inv_2
X_14559_ _25104_/Q _14075_/X _14069_/X VGND VGND VPWR VPWR _14559_/X sky130_fd_sc_hd__a21bo_4
XFILLER_159_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17278_ _17203_/Y _17243_/X _17277_/X VGND VGND VPWR VPWR _17278_/X sky130_fd_sc_hd__or3_4
XFILLER_147_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23038__A2 _22851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_121_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24073_/CLK sky130_fd_sc_hd__clkbuf_1
X_16229_ _16229_/A VGND VGND VPWR VPWR _16229_/Y sky130_fd_sc_hd__inv_2
X_19017_ _23896_/Q VGND VGND VPWR VPWR _19017_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_184_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _25491_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22797__B2 _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19919_ _19919_/A VGND VGND VPWR VPWR _21495_/B sky130_fd_sc_hd__inv_2
XFILLER_96_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22930_ _22930_/A _22928_/X _22929_/X VGND VGND VPWR VPWR _22930_/X sky130_fd_sc_hd__or3_4
XANTENNA__14239__B1 _13849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22861_ _21719_/B VGND VGND VPWR VPWR _22861_/X sky130_fd_sc_hd__buf_2
XANTENNA__15987__B1 _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24838__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24600_ _24601_/CLK _16426_/X HRESETn VGND VGND VPWR VPWR _24600_/Q sky130_fd_sc_hd__dfrtp_4
X_21812_ _21482_/A _21812_/B _21811_/X VGND VGND VPWR VPWR _21812_/X sky130_fd_sc_hd__and3_4
X_22792_ _22792_/A _22662_/B VGND VGND VPWR VPWR _22792_/X sky130_fd_sc_hd__or2_4
XFILLER_225_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17728__B2 _21675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24531_ _24566_/CLK _24531_/D HRESETn VGND VGND VPWR VPWR _16603_/A sky130_fd_sc_hd__dfrtp_4
X_21743_ _18388_/Y _12080_/X _12125_/Y _21579_/X VGND VGND VPWR VPWR _21743_/X sky130_fd_sc_hd__o22a_4
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22684__B _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24462_ _25023_/CLK _24462_/D HRESETn VGND VGND VPWR VPWR _24462_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21674_ _21482_/A _21672_/X _21674_/C VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__and3_4
XFILLER_12_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23590_/CLK _23413_/D VGND VGND VPWR VPWR _20379_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20625_ _14877_/Y _20623_/X _20680_/A _20624_/X VGND VGND VPWR VPWR _20626_/A sky130_fd_sc_hd__a211o_4
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24393_ _24406_/CLK _17124_/X HRESETn VGND VGND VPWR VPWR _24393_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23344_ _23253_/A _23341_/X _23344_/C VGND VGND VPWR VPWR _23349_/C sky130_fd_sc_hd__and3_4
X_20556_ _18891_/X VGND VGND VPWR VPWR _20556_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_80_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_80_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23275_ _24480_/Q _22968_/B _22853_/X VGND VGND VPWR VPWR _23275_/X sky130_fd_sc_hd__and3_4
XANTENNA__15911__B1 _15632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20487_ _20487_/A _20487_/B VGND VGND VPWR VPWR _20533_/C sky130_fd_sc_hd__or2_4
X_25014_ _25011_/CLK _25014_/D HRESETn VGND VGND VPWR VPWR _25014_/Q sky130_fd_sc_hd__dfrtp_4
X_22226_ _22226_/A _18919_/Y VGND VGND VPWR VPWR _22226_/X sky130_fd_sc_hd__or2_4
XANTENNA__22205__A _22171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22157_ _22146_/B _22155_/X _22157_/C VGND VGND VPWR VPWR _22157_/X sky130_fd_sc_hd__and3_4
XFILLER_105_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21108_ _21747_/A _21107_/Y _24649_/Q _21747_/A VGND VGND VPWR VPWR _21108_/X sky130_fd_sc_hd__a2bb2o_4
X_22088_ _21257_/A VGND VGND VPWR VPWR _22385_/A sky130_fd_sc_hd__buf_2
XFILLER_219_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13930_ _24980_/Q VGND VGND VPWR VPWR _13964_/A sky130_fd_sc_hd__inv_2
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21039_ _22541_/A VGND VGND VPWR VPWR _21039_/X sky130_fd_sc_hd__buf_2
XFILLER_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13861_ _24007_/Q VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__buf_2
XFILLER_247_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23036__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24579__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15600_ _22934_/A _15597_/X _11793_/X _15597_/X VGND VGND VPWR VPWR _15600_/X sky130_fd_sc_hd__a2bb2o_4
X_12812_ _12912_/B _22726_/A _12912_/B _22726_/A VGND VGND VPWR VPWR _12813_/D sky130_fd_sc_hd__a2bb2o_4
X_16580_ _16578_/Y _16579_/X _16410_/X _16579_/X VGND VGND VPWR VPWR _24541_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ _13792_/A VGND VGND VPWR VPWR _13793_/D sky130_fd_sc_hd__buf_2
XFILLER_43_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ _15530_/Y _15526_/X HADDR[10] _15526_/X VGND VGND VPWR VPWR _15531_/X sky130_fd_sc_hd__a2bb2o_4
X_12743_ _12740_/B _12742_/Y _12741_/C VGND VGND VPWR VPWR _12743_/X sky130_fd_sc_hd__and3_4
X_24729_ _24732_/CLK _24729_/D HRESETn VGND VGND VPWR VPWR _24729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18250_ _11706_/Y _18243_/X _15756_/X _18243_/X VGND VGND VPWR VPWR _24244_/D sky130_fd_sc_hd__a2bb2o_4
X_15462_ _13955_/A _15458_/X _15455_/X _13963_/B _15461_/X VGND VGND VPWR VPWR _24970_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _12710_/B _12627_/X VGND VGND VPWR VPWR _12674_/X sky130_fd_sc_hd__or2_4
XANTENNA__23268__A2 _21890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _24365_/Q VGND VGND VPWR VPWR _17263_/C sky130_fd_sc_hd__inv_2
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _20610_/A _14392_/X _14412_/X _14392_/X VGND VGND VPWR VPWR _14413_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18181_ _17977_/A _18181_/B VGND VGND VPWR VPWR _18181_/X sky130_fd_sc_hd__or2_4
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15393_/A _15391_/X _15392_/X VGND VGND VPWR VPWR _24994_/D sky130_fd_sc_hd__and3_4
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _17132_/A _17132_/B VGND VGND VPWR VPWR _17133_/C sky130_fd_sc_hd__or2_4
XFILLER_129_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _25172_/Q _14342_/X VGND VGND VPWR VPWR _14349_/D sky130_fd_sc_hd__or2_4
XANTENNA__25146__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16155__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063_ _17095_/A _17061_/X _17062_/Y VGND VGND VPWR VPWR _24409_/D sky130_fd_sc_hd__and3_4
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14275_ _25194_/Q VGND VGND VPWR VPWR _14275_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16014_ _24749_/Q VGND VGND VPWR VPWR _16014_/Y sky130_fd_sc_hd__inv_2
X_13226_ _13423_/A VGND VGND VPWR VPWR _13391_/A sky130_fd_sc_hd__buf_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15936__B _15934_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13157_ _13178_/A VGND VGND VPWR VPWR _13195_/A sky130_fd_sc_hd__buf_2
XANTENNA__14469__B1 _14427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12108_ _16193_/A _12108_/B VGND VGND VPWR VPWR _12108_/X sky130_fd_sc_hd__or2_4
X_13088_ _13088_/A _12992_/Y VGND VGND VPWR VPWR _13115_/B sky130_fd_sc_hd__or2_4
X_17965_ _17943_/A _17965_/B VGND VGND VPWR VPWR _17965_/X sky130_fd_sc_hd__or2_4
X_19704_ _19698_/Y VGND VGND VPWR VPWR _19704_/X sky130_fd_sc_hd__buf_2
XANTENNA__15952__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12039_ _11998_/Y _12038_/X _25499_/Q _12038_/X VGND VGND VPWR VPWR _12039_/X sky130_fd_sc_hd__a2bb2o_4
X_16916_ _24271_/Q VGND VGND VPWR VPWR _16916_/Y sky130_fd_sc_hd__inv_2
X_17896_ _17896_/A _17858_/B _17895_/X VGND VGND VPWR VPWR _24263_/D sky130_fd_sc_hd__and3_4
XFILLER_214_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19635_ _23681_/Q VGND VGND VPWR VPWR _19635_/Y sky130_fd_sc_hd__inv_2
X_16847_ _16845_/Y _16846_/X _15761_/X _16846_/X VGND VGND VPWR VPWR _16847_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15969__B1 _15967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ _11865_/X VGND VGND VPWR VPWR _19566_/X sky130_fd_sc_hd__buf_2
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16778_ _24462_/Q VGND VGND VPWR VPWR _16778_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_23_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22703__A1 _12247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18517_ _18517_/A _18517_/B VGND VGND VPWR VPWR _18517_/X sky130_fd_sc_hd__or2_4
XFILLER_240_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15729_ _12591_/Y _15727_/X _11763_/X _15727_/X VGND VGND VPWR VPWR _24888_/D sky130_fd_sc_hd__a2bb2o_4
X_19497_ _21691_/B _19496_/X _11961_/X _19496_/X VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18448_ _16209_/Y _24189_/Q _16224_/A _18531_/A VGND VGND VPWR VPWR _18451_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16394__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12404__C1 _12403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18379_ _18379_/A VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__buf_2
XANTENNA__14944__B2 _14943_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19332__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20410_ _23401_/Q VGND VGND VPWR VPWR _20410_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21390_ _21248_/A VGND VGND VPWR VPWR _21408_/A sky130_fd_sc_hd__buf_2
XANTENNA__16146__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22951__C _22944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20341_ _20340_/Y _20336_/X _20034_/X _20323_/Y VGND VGND VPWR VPWR _20341_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20272_ _13414_/B VGND VGND VPWR VPWR _20272_/Y sky130_fd_sc_hd__inv_2
X_23060_ _23060_/A VGND VGND VPWR VPWR _23060_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19852__A2_N _19851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22011_ _13793_/D _23358_/B VGND VGND VPWR VPWR _22011_/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16449__B2 _16446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23962_ _25215_/CLK _20608_/Y HRESETn VGND VGND VPWR VPWR _18875_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21583__B _21583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22913_ _22913_/A _22985_/B VGND VGND VPWR VPWR _22913_/X sky130_fd_sc_hd__or2_4
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24672__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23893_ _24101_/CLK _19025_/X VGND VGND VPWR VPWR _19024_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14478__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22844_ _23087_/B VGND VGND VPWR VPWR _22844_/X sky130_fd_sc_hd__buf_2
XANTENNA__24601__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22775_ _22774_/X VGND VGND VPWR VPWR _22775_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22170__A2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19571__B1 _19410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24514_ _24509_/CLK _24514_/D HRESETn VGND VGND VPWR VPWR _16651_/A sky130_fd_sc_hd__dfrtp_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21726_ _21726_/A _21726_/B VGND VGND VPWR VPWR _21730_/A sky130_fd_sc_hd__or2_4
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25494_ _25494_/CLK _25494_/D HRESETn VGND VGND VPWR VPWR _25494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23303__B _23303_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24445_ _24476_/CLK _24445_/D HRESETn VGND VGND VPWR VPWR _24445_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21104__A _24617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21657_ _19614_/A _21971_/B _19564_/A _21656_/X VGND VGND VPWR VPWR _21657_/X sky130_fd_sc_hd__o22a_4
X_20608_ _20608_/A _20608_/B VGND VGND VPWR VPWR _20608_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16137__B1 _11805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12390_ _12390_/A _12390_/B _12380_/X _12389_/X VGND VGND VPWR VPWR _12391_/B sky130_fd_sc_hd__or4_4
X_24376_ _24641_/CLK _24376_/D HRESETn VGND VGND VPWR VPWR _17244_/A sky130_fd_sc_hd__dfrtp_4
X_21588_ _15715_/X VGND VGND VPWR VPWR _21588_/X sky130_fd_sc_hd__buf_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23327_ _23327_/A VGND VGND VPWR VPWR _23327_/Y sky130_fd_sc_hd__inv_2
X_20539_ _24087_/Q _20543_/B _20511_/X VGND VGND VPWR VPWR _20539_/X sky130_fd_sc_hd__a21o_4
XFILLER_165_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14060_ _14060_/A _14060_/B _14060_/C _14059_/X VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__or4_4
X_23258_ _23156_/A _23258_/B _23253_/X _23258_/D VGND VGND VPWR VPWR _23258_/X sky130_fd_sc_hd__or4_4
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13011_ _13011_/A _13021_/C _13010_/X VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__or3_4
X_22209_ _22209_/A _22207_/X _22209_/C VGND VGND VPWR VPWR _22214_/B sky130_fd_sc_hd__and3_4
XFILLER_134_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17029__A _17345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23189_ _24611_/Q _23189_/B VGND VGND VPWR VPWR _23189_/X sky130_fd_sc_hd__or2_4
XANTENNA__12461__A _12247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_24_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _23590_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_87_0_HCLK clkbuf_8_86_0_HCLK/A VGND VGND VPWR VPWR _25358_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_239_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16868__A _14791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22589__B _22589_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14962_ _14962_/A VGND VGND VPWR VPWR _15251_/A sky130_fd_sc_hd__buf_2
X_17750_ _24289_/Q VGND VGND VPWR VPWR _17750_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16701_ _16701_/A VGND VGND VPWR VPWR _22616_/A sky130_fd_sc_hd__inv_2
X_13913_ _13955_/B VGND VGND VPWR VPWR _13913_/Y sky130_fd_sc_hd__inv_2
X_14893_ pwm_S6 VGND VGND VPWR VPWR _14893_/Y sky130_fd_sc_hd__inv_2
X_17681_ _17585_/C _17683_/B _17680_/Y VGND VGND VPWR VPWR _17681_/X sky130_fd_sc_hd__o21a_4
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19420_ _23754_/Q VGND VGND VPWR VPWR _19420_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11805__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13844_ _13844_/A VGND VGND VPWR VPWR _13844_/X sky130_fd_sc_hd__buf_2
X_16632_ _21167_/A _16554_/A _16375_/X _16554_/A VGND VGND VPWR VPWR _16632_/X sky130_fd_sc_hd__a2bb2o_4
X_19351_ _19350_/Y _19348_/X _19305_/X _19348_/X VGND VGND VPWR VPWR _19351_/X sky130_fd_sc_hd__a2bb2o_4
X_13775_ _13760_/X VGND VGND VPWR VPWR _13775_/X sky130_fd_sc_hd__buf_2
X_16563_ _16562_/Y _16560_/X _16393_/X _16560_/X VGND VGND VPWR VPWR _16563_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18302_ _18301_/X VGND VGND VPWR VPWR _18302_/Y sky130_fd_sc_hd__inv_2
XFILLER_215_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ _12728_/A _12723_/B _12726_/C VGND VGND VPWR VPWR _12726_/X sky130_fd_sc_hd__and3_4
X_15514_ _15512_/Y _15508_/X HADDR[17] _15513_/X VGND VGND VPWR VPWR _15514_/X sky130_fd_sc_hd__a2bb2o_4
X_16494_ _24573_/Q VGND VGND VPWR VPWR _16494_/Y sky130_fd_sc_hd__inv_2
X_19282_ _19277_/Y _19281_/X _16872_/X _19281_/X VGND VGND VPWR VPWR _23804_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16376__B1 _16375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15445_ _13958_/A _15441_/X _15444_/X VGND VGND VPWR VPWR _15445_/Y sky130_fd_sc_hd__o21ai_4
X_18233_ _18169_/A _18233_/B _18233_/C VGND VGND VPWR VPWR _18234_/C sky130_fd_sc_hd__and3_4
XANTENNA__25548__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12657_ _12657_/A _12657_/B _12656_/X VGND VGND VPWR VPWR _12658_/A sky130_fd_sc_hd__or3_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14926__B2 _14925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19314__B1 _19246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15376_ _15376_/A _15376_/B VGND VGND VPWR VPWR _15376_/Y sky130_fd_sc_hd__nand2_4
X_18164_ _18164_/A _19158_/A VGND VGND VPWR VPWR _18166_/B sky130_fd_sc_hd__or2_4
XFILLER_191_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12588_ _12588_/A VGND VGND VPWR VPWR _12588_/Y sky130_fd_sc_hd__inv_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _14315_/A _14326_/X _25325_/Q _14320_/X VGND VGND VPWR VPWR _14327_/X sky130_fd_sc_hd__o22a_4
X_17115_ _17118_/A _17115_/B VGND VGND VPWR VPWR _17119_/B sky130_fd_sc_hd__or2_4
X_18095_ _18130_/A _18093_/X _18095_/C VGND VGND VPWR VPWR _18095_/X sky130_fd_sc_hd__and3_4
XFILLER_7_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15947__A _15947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17046_ _24390_/Q VGND VGND VPWR VPWR _17129_/A sky130_fd_sc_hd__inv_2
X_14258_ _23979_/Q _13940_/Y VGND VGND VPWR VPWR _15437_/A sky130_fd_sc_hd__or2_4
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13209_ _13209_/A VGND VGND VPWR VPWR _13209_/X sky130_fd_sc_hd__buf_2
X_14189_ _14188_/X VGND VGND VPWR VPWR _25216_/D sky130_fd_sc_hd__inv_2
X_18997_ _18996_/Y _18992_/X _18908_/X _18992_/X VGND VGND VPWR VPWR _23902_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15682__A _15681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17948_ _17951_/A _23844_/Q VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__or2_4
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17879_ _16920_/Y _17877_/X _17878_/Y VGND VGND VPWR VPWR _17879_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19618_ _21976_/B _19615_/X _19454_/X _19615_/X VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20890_ _20878_/X _20889_/Y _16699_/A _20883_/X VGND VGND VPWR VPWR _20890_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19549_ _21217_/A VGND VGND VPWR VPWR _21382_/B sky130_fd_sc_hd__inv_2
XFILLER_222_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19553__B1 _19439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22560_ _16606_/A _23303_/B _21755_/A _22559_/X VGND VGND VPWR VPWR _22561_/C sky130_fd_sc_hd__a211o_4
XFILLER_179_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21511_ _22400_/A VGND VGND VPWR VPWR _21511_/X sky130_fd_sc_hd__buf_2
XANTENNA__25289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22491_ _22488_/X _22490_/X _21434_/X _24869_/Q _22558_/A VGND VGND VPWR VPWR _22492_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18108__A1 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24230_ _24230_/CLK _24230_/D HRESETn VGND VGND VPWR VPWR _18267_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21442_ _15866_/X VGND VGND VPWR VPWR _21543_/A sky130_fd_sc_hd__buf_2
XANTENNA__16119__B1 _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21112__B1 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24161_ _25212_/CLK _24161_/D HRESETn VGND VGND VPWR VPWR _24161_/Q sky130_fd_sc_hd__dfrtp_4
X_21373_ _21373_/A VGND VGND VPWR VPWR _21733_/B sky130_fd_sc_hd__buf_2
XFILLER_175_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14761__A _14761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23112_ _23089_/X _23112_/B _23112_/C _23111_/X VGND VGND VPWR VPWR HRDATA[24] sky130_fd_sc_hd__or4_4
XFILLER_207_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20324_ _20323_/Y VGND VGND VPWR VPWR _20324_/X sky130_fd_sc_hd__buf_2
X_24092_ _24966_/CLK _24092_/D HRESETn VGND VGND VPWR VPWR _20487_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23043_ _12833_/Y _22725_/X _22291_/B _12595_/Y _22862_/X VGND VGND VPWR VPWR _23043_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_162_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20255_ _20255_/A VGND VGND VPWR VPWR _20255_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_240_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24160_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_88_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20186_ _23486_/Q VGND VGND VPWR VPWR _21407_/B sky130_fd_sc_hd__inv_2
XANTENNA__24853__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16802__A2_N _16738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24994_ _24975_/CLK _24994_/D HRESETn VGND VGND VPWR VPWR _24994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23945_ _23946_/CLK _20991_/X HRESETn VGND VGND VPWR VPWR _20995_/B sky130_fd_sc_hd__dfstp_4
XANTENNA__13824__B _17422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11890_ _11889_/Y VGND VGND VPWR VPWR _11890_/X sky130_fd_sc_hd__buf_2
X_23876_ _24214_/CLK _19078_/X VGND VGND VPWR VPWR _23876_/Q sky130_fd_sc_hd__dfxtp_4
X_22827_ _16231_/A _22827_/B VGND VGND VPWR VPWR _22832_/B sky130_fd_sc_hd__or2_4
XANTENNA__22679__B1 _17762_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13560_ _25266_/Q VGND VGND VPWR VPWR _13560_/Y sky130_fd_sc_hd__inv_2
X_25546_ _24697_/CLK _25546_/D HRESETn VGND VGND VPWR VPWR _25546_/Q sky130_fd_sc_hd__dfrtp_4
X_22758_ _22758_/A _22789_/B VGND VGND VPWR VPWR _22758_/X sky130_fd_sc_hd__or2_4
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12511_ _12232_/Y _12514_/B VGND VGND VPWR VPWR _12512_/C sky130_fd_sc_hd__nand2_4
XFILLER_197_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21709_ _21709_/A _23016_/A VGND VGND VPWR VPWR _21709_/X sky130_fd_sc_hd__or2_4
XFILLER_185_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13491_ _13486_/A VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__buf_2
X_25477_ _24119_/CLK _12126_/X HRESETn VGND VGND VPWR VPWR _12125_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22689_ _16284_/X _22689_/B VGND VGND VPWR VPWR _22689_/Y sky130_fd_sc_hd__nor2_4
XFILLER_157_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15230_ _14935_/X _15228_/X _15229_/Y VGND VGND VPWR VPWR _25032_/D sky130_fd_sc_hd__o21a_4
X_12442_ _12269_/Y _12442_/B VGND VGND VPWR VPWR _12442_/X sky130_fd_sc_hd__or2_4
X_24428_ _25018_/CLK _16850_/X HRESETn VGND VGND VPWR VPWR _24428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19847__B2 _19844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15161_ _15152_/X _15155_/X _15161_/C _15161_/D VGND VGND VPWR VPWR _15161_/X sky130_fd_sc_hd__or4_4
XFILLER_172_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15767__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12373_ _24853_/Q VGND VGND VPWR VPWR _12373_/Y sky130_fd_sc_hd__inv_2
X_24359_ _24346_/CLK _17350_/X HRESETn VGND VGND VPWR VPWR _17348_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_50_0_HCLK clkbuf_6_50_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _14112_/A _14112_/B _25228_/Q VGND VGND VPWR VPWR _14112_/X sky130_fd_sc_hd__or3_4
XFILLER_126_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15092_ _15092_/A VGND VGND VPWR VPWR _15092_/Y sky130_fd_sc_hd__inv_2
X_14043_ _14043_/A _14032_/B _14042_/X _14034_/D VGND VGND VPWR VPWR _14043_/X sky130_fd_sc_hd__or4_4
X_18920_ _18919_/Y _18917_/X _16876_/X _18917_/X VGND VGND VPWR VPWR _18920_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18851_ _18851_/A _18840_/X _18845_/X _18850_/X VGND VGND VPWR VPWR _18851_/X sky130_fd_sc_hd__or4_4
XFILLER_192_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24594__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17802_ _16952_/Y _17770_/X _17562_/X VGND VGND VPWR VPWR _17802_/X sky130_fd_sc_hd__or3_4
XANTENNA__24523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _18782_/A _18782_/B VGND VGND VPWR VPWR _18784_/B sky130_fd_sc_hd__or2_4
XFILLER_209_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15994_ _15797_/X _15895_/A _15993_/X _21715_/A _15940_/X VGND VGND VPWR VPWR _24756_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22112__B _22176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17733_ _17733_/A _17720_/X VGND VGND VPWR VPWR _17733_/X sky130_fd_sc_hd__and2_4
X_14945_ _25015_/Q VGND VGND VPWR VPWR _15290_/A sky130_fd_sc_hd__inv_2
XANTENNA__16942__A1_N _16143_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17664_ _17581_/Y _17664_/B VGND VGND VPWR VPWR _17667_/B sky130_fd_sc_hd__or2_4
XFILLER_235_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14876_ _14820_/X _14875_/Y _24959_/Q _14820_/X VGND VGND VPWR VPWR _14876_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19403_ _19401_/Y _19397_/X _19402_/X _19397_/X VGND VGND VPWR VPWR _19403_/X sky130_fd_sc_hd__a2bb2o_4
X_16615_ _16615_/A VGND VGND VPWR VPWR _16615_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ _13826_/X VGND VGND VPWR VPWR _13828_/D sky130_fd_sc_hd__buf_2
X_17595_ _17566_/Y _17595_/B VGND VGND VPWR VPWR _17596_/B sky130_fd_sc_hd__nor2_4
X_19334_ _19333_/Y _19331_/X _19220_/X _19331_/X VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13758_ _13757_/C VGND VGND VPWR VPWR _18914_/A sky130_fd_sc_hd__inv_2
X_16546_ _24553_/Q VGND VGND VPWR VPWR _16546_/Y sky130_fd_sc_hd__inv_2
X_12709_ _12708_/X VGND VGND VPWR VPWR _12709_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19265_ _22070_/B _19259_/X _16881_/X _19264_/X VGND VGND VPWR VPWR _23810_/D sky130_fd_sc_hd__a2bb2o_4
X_13689_ _13688_/Y VGND VGND VPWR VPWR _13689_/X sky130_fd_sc_hd__buf_2
X_16477_ _16474_/Y _16470_/X _16389_/X _16476_/X VGND VGND VPWR VPWR _16477_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18216_ _17984_/A _19477_/A VGND VGND VPWR VPWR _18216_/X sky130_fd_sc_hd__or2_4
XANTENNA__25311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15428_ _15424_/A _15424_/B VGND VGND VPWR VPWR _15429_/B sky130_fd_sc_hd__nand2_4
XANTENNA__21679__A _21679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19196_ _19196_/A VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__buf_2
XFILLER_163_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15359_ _15387_/A VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__buf_2
X_18147_ _17988_/A _18145_/X _18146_/X VGND VGND VPWR VPWR _18148_/C sky130_fd_sc_hd__and3_4
XFILLER_144_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25202__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18078_ _17988_/A _18078_/B _18077_/X VGND VGND VPWR VPWR _18078_/X sky130_fd_sc_hd__and3_4
XANTENNA__16521__B1 _16252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17029_ _17345_/A VGND VGND VPWR VPWR _17064_/A sky130_fd_sc_hd__buf_2
XFILLER_236_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20040_ _22347_/B _20039_/X _19990_/X _20039_/X VGND VGND VPWR VPWR _23540_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18274__B1 _16861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_70_0_HCLK clkbuf_8_70_0_HCLK/A VGND VGND VPWR VPWR _24777_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13644__B _14679_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21991_ _18357_/A _21991_/B VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__and2_4
XANTENNA__22957__B _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19774__B1 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23730_ _23441_/CLK _19490_/X VGND VGND VPWR VPWR _19488_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _20927_/X _20941_/Y _16669_/A _20931_/X VGND VGND VPWR VPWR _24071_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_215_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19612__A _11861_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23642_/CLK _19695_/X VGND VGND VPWR VPWR _13457_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_198_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20872_/X VGND VGND VPWR VPWR _24055_/D sky130_fd_sc_hd__inv_2
XFILLER_199_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25400_ _25402_/CLK _25400_/D HRESETn VGND VGND VPWR VPWR _12888_/A sky130_fd_sc_hd__dfrtp_4
X_22612_ _21082_/A _22609_/X _21116_/X _22611_/X VGND VGND VPWR VPWR _22612_/Y sky130_fd_sc_hd__a22oi_4
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23560_/CLK _23592_/D VGND VGND VPWR VPWR _23592_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25331_ _25507_/CLK _13473_/X HRESETn VGND VGND VPWR VPWR _25331_/Q sky130_fd_sc_hd__dfrtp_4
X_22543_ _22543_/A VGND VGND VPWR VPWR _22543_/X sky130_fd_sc_hd__buf_2
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25262_ _25276_/CLK _25262_/D HRESETn VGND VGND VPWR VPWR _25262_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21589__A _15019_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22474_ _21605_/A VGND VGND VPWR VPWR _23144_/A sky130_fd_sc_hd__buf_2
XANTENNA__16760__B1 _16412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24213_ _23459_/CLK _24213_/D HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _21338_/X _21425_/B _21425_/C _21425_/D VGND VGND VPWR VPWR _21425_/X sky130_fd_sc_hd__or4_4
X_25193_ _25253_/CLK _25193_/D HRESETn VGND VGND VPWR VPWR _14277_/A sky130_fd_sc_hd__dfrtp_4
X_24144_ _24145_/CLK _24144_/D HRESETn VGND VGND VPWR VPWR _18782_/A sky130_fd_sc_hd__dfrtp_4
X_21356_ _14229_/A VGND VGND VPWR VPWR _21356_/X sky130_fd_sc_hd__buf_2
XFILLER_146_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20307_ _23441_/Q VGND VGND VPWR VPWR _20307_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24075_ _24073_/CLK _20959_/X HRESETn VGND VGND VPWR VPWR _20956_/A sky130_fd_sc_hd__dfrtp_4
X_21287_ _13607_/B VGND VGND VPWR VPWR _22523_/A sky130_fd_sc_hd__buf_2
X_23026_ _17231_/A _21065_/X VGND VGND VPWR VPWR _23029_/B sky130_fd_sc_hd__or2_4
XANTENNA__18265__B1 _16726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23300__A2_N _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20238_ _20237_/Y _20235_/X _19769_/X _20235_/X VGND VGND VPWR VPWR _23467_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20169_ _20169_/A VGND VGND VPWR VPWR _20169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18280__A3 _13481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12991_ _13051_/A VGND VGND VPWR VPWR _13044_/A sky130_fd_sc_hd__buf_2
X_24977_ _24979_/CLK _15451_/X HRESETn VGND VGND VPWR VPWR _13942_/A sky130_fd_sc_hd__dfrtp_4
X_11942_ _19632_/A VGND VGND VPWR VPWR _11942_/Y sky130_fd_sc_hd__inv_2
X_14730_ _13753_/X _14713_/Y _14730_/C VGND VGND VPWR VPWR _14730_/X sky130_fd_sc_hd__and3_4
XFILLER_85_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23928_ _23577_/CLK _18927_/X VGND VGND VPWR VPWR _18926_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_233_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14661_ _17944_/A VGND VGND VPWR VPWR _17951_/A sky130_fd_sc_hd__buf_2
X_11873_ _25525_/Q VGND VGND VPWR VPWR _11873_/Y sky130_fd_sc_hd__inv_2
X_23859_ _24111_/CLK _23859_/D VGND VGND VPWR VPWR _13215_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13612_ _25080_/Q VGND VGND VPWR VPWR _13613_/B sky130_fd_sc_hd__buf_2
X_16400_ _24610_/Q VGND VGND VPWR VPWR _16400_/Y sky130_fd_sc_hd__inv_2
X_14592_ _14590_/X _14566_/X _14591_/X _13779_/X _14586_/C VGND VGND VPWR VPWR _25101_/D
+ sky130_fd_sc_hd__a32o_4
X_17380_ _17380_/A VGND VGND VPWR VPWR _17380_/Y sky130_fd_sc_hd__inv_2
X_13543_ _13543_/A VGND VGND VPWR VPWR _13543_/Y sky130_fd_sc_hd__inv_2
X_16331_ _24633_/Q VGND VGND VPWR VPWR _16331_/Y sky130_fd_sc_hd__inv_2
X_25529_ _25528_/CLK _25529_/D HRESETn VGND VGND VPWR VPWR _11853_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16262_ _16261_/Y _16257_/X _16066_/X _16257_/X VGND VGND VPWR VPWR _24659_/D sky130_fd_sc_hd__a2bb2o_4
X_19050_ _19050_/A VGND VGND VPWR VPWR _19050_/Y sky130_fd_sc_hd__inv_2
X_13474_ _13474_/A VGND VGND VPWR VPWR _13474_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23077__B1 _22816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16751__B1 _15734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22419__A3 _22148_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15213_ _15068_/X _15202_/X _15213_/C VGND VGND VPWR VPWR _25036_/D sky130_fd_sc_hd__and3_4
X_18001_ _18158_/A _23907_/Q VGND VGND VPWR VPWR _18002_/C sky130_fd_sc_hd__or2_4
X_12425_ _12425_/A _12425_/B VGND VGND VPWR VPWR _12428_/B sky130_fd_sc_hd__or2_4
XANTENNA__12368__B2 _24840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16193_ _16193_/A _22462_/A VGND VGND VPWR VPWR _16193_/X sky130_fd_sc_hd__or2_4
XFILLER_138_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12914__A _12834_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15144_ _15354_/A VGND VGND VPWR VPWR _15346_/A sky130_fd_sc_hd__inv_2
X_12356_ _12356_/A VGND VGND VPWR VPWR _13006_/B sky130_fd_sc_hd__inv_2
XFILLER_154_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16503__B1 _16417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24775__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15857__A2 _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15075_ _14969_/Y _14958_/Y _15075_/C _15075_/D VGND VGND VPWR VPWR _15075_/X sky130_fd_sc_hd__or4_4
X_19952_ _19950_/Y _19946_/X _19632_/X _19951_/X VGND VGND VPWR VPWR _19952_/X sky130_fd_sc_hd__a2bb2o_4
X_12287_ _12287_/A _12238_/Y _12263_/Y _12205_/Y VGND VGND VPWR VPWR _12287_/X sky130_fd_sc_hd__or4_4
XANTENNA__24704__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14026_ _14033_/A VGND VGND VPWR VPWR _14026_/Y sky130_fd_sc_hd__inv_2
X_18903_ _18901_/Y _18902_/Y _17452_/X _18902_/Y VGND VGND VPWR VPWR _24122_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22052__A1 _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18256__B1 _16613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19883_ _19895_/A VGND VGND VPWR VPWR _19883_/X sky130_fd_sc_hd__buf_2
XFILLER_141_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22052__B2 _22051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18834_ _16478_/Y _24159_/Q _16478_/Y _24159_/Q VGND VGND VPWR VPWR _18834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_57_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18765_ _18765_/A _18769_/B VGND VGND VPWR VPWR _18765_/Y sky130_fd_sc_hd__nand2_4
X_15977_ _15863_/X VGND VGND VPWR VPWR _15977_/X sky130_fd_sc_hd__buf_2
XANTENNA__15490__B1 _15489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17716_ _17716_/A VGND VGND VPWR VPWR _21485_/A sky130_fd_sc_hd__buf_2
XANTENNA__15960__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14928_ _24443_/Q VGND VGND VPWR VPWR _14928_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18696_ _18694_/Y _18772_/A _18617_/Y _18696_/D VGND VGND VPWR VPWR _18699_/C sky130_fd_sc_hd__or4_4
XFILLER_48_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17647_ _17516_/Y _17652_/B _17600_/X VGND VGND VPWR VPWR _17647_/Y sky130_fd_sc_hd__a21oi_4
X_14859_ _14837_/X _14858_/X _25199_/Q _14844_/X VGND VGND VPWR VPWR _14859_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17578_ _17531_/Y _17578_/B _17577_/X VGND VGND VPWR VPWR _17579_/C sky130_fd_sc_hd__or3_4
XANTENNA__22793__A _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19317_ _19315_/Y _19316_/X _19226_/X _19316_/X VGND VGND VPWR VPWR _19317_/X sky130_fd_sc_hd__a2bb2o_4
X_16529_ _16529_/A VGND VGND VPWR VPWR _16529_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17887__A _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16791__A _19085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19248_ _13381_/B VGND VGND VPWR VPWR _19248_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12359__B2 _24839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19179_ _19178_/Y _19174_/X _19131_/X _19174_/X VGND VGND VPWR VPWR _23840_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21210_ _21210_/A _21210_/B VGND VGND VPWR VPWR _21212_/B sky130_fd_sc_hd__or2_4
X_22190_ _25255_/Q _22190_/B VGND VGND VPWR VPWR _22190_/X sky130_fd_sc_hd__and2_4
X_21141_ _14439_/Y _14229_/A _21139_/Y _21353_/A VGND VGND VPWR VPWR _21141_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21072_ _24719_/Q _15662_/Y _21049_/X _21071_/X VGND VGND VPWR VPWR _21073_/A sky130_fd_sc_hd__a211o_4
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23129__A _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22033__A _22029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20023_ _20021_/Y _20017_/X _19996_/X _20022_/X VGND VGND VPWR VPWR _20023_/X sky130_fd_sc_hd__a2bb2o_4
X_24900_ _24485_/CLK _15644_/X HRESETn VGND VGND VPWR VPWR _15643_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17127__A _17064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12531__B2 _24876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24831_ _24849_/CLK _24831_/D HRESETn VGND VGND VPWR VPWR _24831_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15481__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15870__A _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24762_ _24759_/CLK _24762_/D HRESETn VGND VGND VPWR VPWR _22483_/A sky130_fd_sc_hd__dfrtp_4
X_21974_ _21974_/A _21974_/B VGND VGND VPWR VPWR _21974_/Y sky130_fd_sc_hd__nand2_4
XFILLER_227_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23713_ _23408_/CLK _23713_/D VGND VGND VPWR VPWR _23713_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_227_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _24067_/Q _20918_/X _20924_/X VGND VGND VPWR VPWR _20925_/Y sky130_fd_sc_hd__a21oi_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24693_ _24732_/CLK _24693_/D HRESETn VGND VGND VPWR VPWR _22413_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ _23644_/CLK _19744_/X VGND VGND VPWR VPWR _13175_/B sky130_fd_sc_hd__dfxtp_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20856_ _20855_/Y _20850_/Y _13667_/B VGND VGND VPWR VPWR _20856_/X sky130_fd_sc_hd__o21a_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23494_/CLK _23575_/D VGND VGND VPWR VPWR _23575_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20787_ _20761_/X _20786_/Y _24918_/Q _20765_/X VGND VGND VPWR VPWR _20787_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25314_ _24196_/CLK _13522_/X HRESETn VGND VGND VPWR VPWR _13520_/A sky130_fd_sc_hd__dfrtp_4
X_22526_ _22523_/X _22524_/X _21968_/A _22525_/Y VGND VGND VPWR VPWR _22529_/A sky130_fd_sc_hd__o22a_4
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15536__B2 _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25245_ _24340_/CLK _14077_/X HRESETn VGND VGND VPWR VPWR _25245_/Q sky130_fd_sc_hd__dfrtp_4
X_22457_ _21324_/X VGND VGND VPWR VPWR _22510_/C sky130_fd_sc_hd__buf_2
XFILLER_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _12208_/A _22871_/A _12208_/Y _12209_/Y VGND VGND VPWR VPWR _12210_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17289__A1 _17243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21408_ _21408_/A _19940_/Y VGND VGND VPWR VPWR _21409_/C sky130_fd_sc_hd__or2_4
X_13190_ _13177_/A _13188_/X _13189_/X VGND VGND VPWR VPWR _13190_/X sky130_fd_sc_hd__and3_4
X_25176_ _25177_/CLK _25176_/D HRESETn VGND VGND VPWR VPWR _25176_/Q sky130_fd_sc_hd__dfrtp_4
X_22388_ _22388_/A _20148_/Y VGND VGND VPWR VPWR _22390_/B sky130_fd_sc_hd__or2_4
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12141_ _12135_/B VGND VGND VPWR VPWR _12141_/Y sky130_fd_sc_hd__inv_2
X_24127_ _23946_/CLK _18896_/X HRESETn VGND VGND VPWR VPWR _24127_/Q sky130_fd_sc_hd__dfstp_4
X_21339_ _21874_/A VGND VGND VPWR VPWR _22316_/B sky130_fd_sc_hd__buf_2
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12072_ _12072_/A VGND VGND VPWR VPWR _12072_/Y sky130_fd_sc_hd__inv_2
X_24058_ _24532_/CLK _20887_/X HRESETn VGND VGND VPWR VPWR _13670_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23039__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15900_ _15894_/X _15895_/X _16245_/A _22669_/A _15896_/X VGND VGND VPWR VPWR _15900_/X
+ sky130_fd_sc_hd__a32o_4
X_23009_ _23009_/A VGND VGND VPWR VPWR _23013_/A sky130_fd_sc_hd__buf_2
XANTENNA__22585__A2 _22678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16880_ _19800_/A VGND VGND VPWR VPWR _16880_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21793__B1 _14758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22878__A _24635_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15831_ _15825_/X _15828_/X _16245_/A _24838_/Q _15826_/X VGND VGND VPWR VPWR _15831_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21782__A _22388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18550_ _18550_/A _18550_/B _18549_/Y VGND VGND VPWR VPWR _24179_/D sky130_fd_sc_hd__and3_4
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12974_ _12952_/D VGND VGND VPWR VPWR _12974_/Y sky130_fd_sc_hd__inv_2
X_15762_ _15758_/X _15751_/X _15761_/X _24871_/Q _15719_/X VGND VGND VPWR VPWR _24871_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20398__A _20385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21545__B1 _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17501_ _17500_/X VGND VGND VPWR VPWR _24328_/D sky130_fd_sc_hd__inv_2
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14713_ _14713_/A VGND VGND VPWR VPWR _14713_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17213__B2 _24351_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11925_ _25516_/Q _11920_/Y VGND VGND VPWR VPWR _11929_/A sky130_fd_sc_hd__and2_4
X_18481_ _24163_/Q VGND VGND VPWR VPWR _18565_/B sky130_fd_sc_hd__inv_2
XFILLER_61_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21888__A1_N _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15693_ _15693_/A VGND VGND VPWR VPWR _15701_/B sky130_fd_sc_hd__inv_2
XFILLER_205_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17432_ _17432_/A VGND VGND VPWR VPWR _17432_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11813__A _16241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11856_ _14400_/A VGND VGND VPWR VPWR _11856_/X sky130_fd_sc_hd__buf_2
X_14644_ _14643_/Y _14631_/Y _14626_/A _14630_/X VGND VGND VPWR VPWR _14644_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _14605_/A _14574_/X VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__or2_4
X_17363_ _17363_/A _17363_/B _17362_/X VGND VGND VPWR VPWR _17363_/X sky130_fd_sc_hd__and3_4
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ HWDATA[21] VGND VGND VPWR VPWR _11787_/X sky130_fd_sc_hd__buf_2
XFILLER_14_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19102_ _19102_/A VGND VGND VPWR VPWR _19102_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16314_ _16314_/A VGND VGND VPWR VPWR _16314_/Y sky130_fd_sc_hd__inv_2
X_13526_ _25312_/Q VGND VGND VPWR VPWR _13526_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17294_ _17294_/A _17294_/B VGND VGND VPWR VPWR _17295_/C sky130_fd_sc_hd__or2_4
XANTENNA__16724__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19033_ _19026_/Y _19030_/X _19032_/X _19030_/X VGND VGND VPWR VPWR _23892_/D sky130_fd_sc_hd__a2bb2o_4
X_13457_ _13356_/A _13457_/B VGND VGND VPWR VPWR _13459_/B sky130_fd_sc_hd__or2_4
X_16245_ _16245_/A VGND VGND VPWR VPWR _16245_/X sky130_fd_sc_hd__buf_2
X_12408_ _25467_/Q _12408_/B VGND VGND VPWR VPWR _12410_/B sky130_fd_sc_hd__or2_4
X_13388_ _13420_/A _23919_/Q VGND VGND VPWR VPWR _13390_/B sky130_fd_sc_hd__or2_4
X_16176_ _16175_/Y _16097_/X _15489_/X _16097_/X VGND VGND VPWR VPWR _16176_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_20_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12339_ _25349_/Q VGND VGND VPWR VPWR _12339_/Y sky130_fd_sc_hd__inv_2
X_15127_ _24603_/Q VGND VGND VPWR VPWR _15127_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15058_ _15178_/A _24482_/Q _15178_/A _24482_/Q VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__a2bb2o_4
X_19935_ _23576_/Q VGND VGND VPWR VPWR _21780_/B sky130_fd_sc_hd__inv_2
XFILLER_141_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14009_ _25245_/Q VGND VGND VPWR VPWR _14058_/C sky130_fd_sc_hd__buf_2
XFILLER_229_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19866_ _23602_/Q VGND VGND VPWR VPWR _19866_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22788__A _22721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18817_ _18806_/A _18810_/B _18816_/X VGND VGND VPWR VPWR _18817_/X sky130_fd_sc_hd__and3_4
X_19797_ _19788_/Y VGND VGND VPWR VPWR _19797_/X sky130_fd_sc_hd__buf_2
XFILLER_209_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19729__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18748_ _18748_/A VGND VGND VPWR VPWR _18748_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_144_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _25276_/CLK sky130_fd_sc_hd__clkbuf_1
X_18679_ _24157_/Q VGND VGND VPWR VPWR _18702_/A sky130_fd_sc_hd__inv_2
XFILLER_24_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20710_ _21757_/A _20695_/X _20704_/X _20709_/X VGND VGND VPWR VPWR _20711_/A sky130_fd_sc_hd__o22a_4
XANTENNA__11723__A _24079_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21690_ _21684_/X _21689_/X _21499_/X VGND VGND VPWR VPWR _21690_/X sky130_fd_sc_hd__o21a_4
XFILLER_196_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20641_ _20640_/X VGND VGND VPWR VPWR _20641_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22954__C _22954_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23360_ _23360_/A _23360_/B VGND VGND VPWR VPWR _23360_/X sky130_fd_sc_hd__and2_4
X_20572_ _14448_/Y _20551_/X _20565_/X _20571_/X VGND VGND VPWR VPWR _20573_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24697__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22311_ _22205_/X _22281_/Y _22311_/C _22310_/X VGND VGND VPWR VPWR HRDATA[6] sky130_fd_sc_hd__or4_4
XFILLER_177_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23291_ _21881_/X _23290_/X _22484_/X _24890_/Q _23120_/X VGND VGND VPWR VPWR _23292_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24626__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22970__B _22967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25030_ _25030_/CLK _25030_/D HRESETn VGND VGND VPWR VPWR _25030_/Q sky130_fd_sc_hd__dfrtp_4
X_22242_ _21278_/X _22222_/X _22237_/X _22240_/Y _22241_/X VGND VGND VPWR VPWR _22242_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20275__B1 _15656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15865__A _15895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12752__B2 _22605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22173_ _16532_/A _21312_/B _21344_/X VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__o21a_4
XFILLER_191_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16158__A1_N _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21124_ _21123_/X VGND VGND VPWR VPWR _21124_/X sky130_fd_sc_hd__buf_2
XFILLER_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21055_ _21046_/X VGND VGND VPWR VPWR _21109_/B sky130_fd_sc_hd__inv_2
XFILLER_247_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20006_ _19988_/Y VGND VGND VPWR VPWR _20006_/X sky130_fd_sc_hd__buf_2
XFILLER_247_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_40_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_40_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24814_ _24812_/CLK _15884_/X HRESETn VGND VGND VPWR VPWR _24814_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21957_ _21472_/A _21957_/B _21957_/C VGND VGND VPWR VPWR _21957_/X sky130_fd_sc_hd__and3_4
X_24745_ _24372_/CLK _16025_/X HRESETn VGND VGND VPWR VPWR _24745_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A _11710_/B _11889_/A VGND VGND VPWR VPWR _11979_/B sky130_fd_sc_hd__or3_4
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20906_/Y _20911_/B _20907_/X VGND VGND VPWR VPWR _20908_/X sky130_fd_sc_hd__o21a_4
X_12690_ _12619_/A _12689_/X VGND VGND VPWR VPWR _12690_/Y sky130_fd_sc_hd__nand2_4
X_24676_ _24674_/CLK _16216_/X HRESETn VGND VGND VPWR VPWR _16214_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _22443_/A _21886_/X _21449_/A _21887_/X VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23628_/CLK _23627_/D VGND VGND VPWR VPWR _23627_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _24048_/Q _24047_/Q _13662_/B VGND VGND VPWR VPWR _20839_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14360_/A VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__buf_2
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23558_ _24937_/CLK _19982_/X VGND VGND VPWR VPWR _23558_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13228_/A VGND VGND VPWR VPWR _13413_/A sky130_fd_sc_hd__buf_2
XFILLER_10_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _17364_/A _22442_/A _12793_/A _22306_/X VGND VGND VPWR VPWR _22509_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _23978_/Q VGND VGND VPWR VPWR _14291_/X sky130_fd_sc_hd__buf_2
XANTENNA__24367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23488_/CLK _23489_/D VGND VGND VPWR VPWR _23489_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13242_ _13153_/X VGND VGND VPWR VPWR _13242_/X sky130_fd_sc_hd__buf_2
X_16030_ _24742_/Q VGND VGND VPWR VPWR _16030_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25228_ _23395_/CLK _14143_/X HRESETn VGND VGND VPWR VPWR _25228_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21777__A _14709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20681__A _20681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20266__B1 _20243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ _13195_/A _13173_/B VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__or2_4
X_25159_ _25168_/CLK _25159_/D HRESETn VGND VGND VPWR VPWR _25159_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15775__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18151__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12124_ _12122_/Y _12123_/X _11856_/X _12123_/X VGND VGND VPWR VPWR _12124_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17981_ _18097_/A VGND VGND VPWR VPWR _17988_/A sky130_fd_sc_hd__buf_2
XANTENNA__12911__B _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19720_ _19719_/Y VGND VGND VPWR VPWR _19720_/X sky130_fd_sc_hd__buf_2
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19959__B1 _19643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12055_ _12055_/A VGND VGND VPWR VPWR _12055_/Y sky130_fd_sc_hd__inv_2
X_16932_ _16932_/A _16932_/B _16922_/X _16931_/X VGND VGND VPWR VPWR _16962_/A sky130_fd_sc_hd__or4_4
XANTENNA__11808__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19651_ _24213_/Q _18342_/A _17463_/X _20256_/D VGND VGND VPWR VPWR _19652_/A sky130_fd_sc_hd__or4_4
XFILLER_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16863_ _14953_/Y _16805_/X _16726_/X _16805_/X VGND VGND VPWR VPWR _24420_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25106__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18602_ _18565_/B _18503_/X _18505_/X _18599_/Y VGND VGND VPWR VPWR _18603_/A sky130_fd_sc_hd__a211o_4
X_15814_ _15790_/X _15804_/X _15734_/X _24850_/Q _15802_/X VGND VGND VPWR VPWR _24850_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19582_ _19582_/A VGND VGND VPWR VPWR _21962_/B sky130_fd_sc_hd__inv_2
XFILLER_203_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16794_ _24454_/Q VGND VGND VPWR VPWR _16794_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19187__B2 _19181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18533_ _24184_/Q _18533_/B VGND VGND VPWR VPWR _18533_/X sky130_fd_sc_hd__or2_4
XFILLER_46_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15745_ _12542_/Y _15741_/X _11793_/X _15744_/X VGND VGND VPWR VPWR _15745_/X sky130_fd_sc_hd__a2bb2o_4
X_12957_ _12984_/A _12957_/B _12957_/C VGND VGND VPWR VPWR _25384_/D sky130_fd_sc_hd__and3_4
XANTENNA__22191__B1 _14235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_217_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24592_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11908_ _17711_/D VGND VGND VPWR VPWR _11908_/Y sky130_fd_sc_hd__inv_2
X_18464_ _24189_/Q VGND VGND VPWR VPWR _18487_/A sky130_fd_sc_hd__inv_2
X_15676_ _15676_/A VGND VGND VPWR VPWR _15676_/X sky130_fd_sc_hd__buf_2
XFILLER_45_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16945__B1 _16138_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18862__A1_N _16532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12888_ _12888_/A _12888_/B VGND VGND VPWR VPWR _12890_/B sky130_fd_sc_hd__or2_4
XPHY_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17396_/X _17410_/X _24343_/Q _24344_/Q _17413_/X VGND VGND VPWR VPWR _24344_/D
+ sky130_fd_sc_hd__a32o_4
X_14627_ _14624_/Y _13647_/X _14626_/Y VGND VGND VPWR VPWR _14639_/B sky130_fd_sc_hd__o21ai_4
XFILLER_221_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11839_ _11837_/Y _11835_/X _11838_/X _11835_/X VGND VGND VPWR VPWR _11839_/X sky130_fd_sc_hd__a2bb2o_4
X_18395_ _24121_/Q _18377_/X _24196_/Q _18391_/X VGND VGND VPWR VPWR _24196_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18326__A _17710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22509__A1_N _17364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17346_ _17258_/Y _17345_/X VGND VGND VPWR VPWR _17347_/A sky130_fd_sc_hd__or2_4
XFILLER_202_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14558_ _14551_/X _14557_/Y sda_oen_o_S4 _14551_/X VGND VGND VPWR VPWR _14558_/X
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24790__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13509_ _12023_/Y _13507_/X _11838_/X _13507_/X VGND VGND VPWR VPWR _13509_/X sky130_fd_sc_hd__a2bb2o_4
X_17277_ _17277_/A _17276_/X VGND VGND VPWR VPWR _17277_/X sky130_fd_sc_hd__or2_4
X_14489_ _25124_/Q VGND VGND VPWR VPWR _14489_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19016_ _19015_/Y _19013_/X _18969_/X _19013_/X VGND VGND VPWR VPWR _23897_/D sky130_fd_sc_hd__a2bb2o_4
X_16228_ _16226_/Y _16222_/X _15967_/X _16227_/X VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21687__A _21687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16159_ _22413_/A VGND VGND VPWR VPWR _16159_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18061__A _18008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18870__B1 _24572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19918_ _19916_/Y _19917_/X _19643_/X _19917_/X VGND VGND VPWR VPWR _23583_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12498__B1 _12403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19849_ _21763_/B _19844_/X _19803_/X _19844_/X VGND VGND VPWR VPWR _19849_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22311__A _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22860_ _23106_/A _22859_/X VGND VGND VPWR VPWR _22860_/Y sky130_fd_sc_hd__nor2_4
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21811_ _21673_/A _21811_/B VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__or2_4
X_22791_ _22791_/A VGND VGND VPWR VPWR _22791_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24530_ _24566_/CLK _24530_/D HRESETn VGND VGND VPWR VPWR _16606_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18925__B2 _18922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21742_ _13518_/Y _21579_/X _12047_/Y _21580_/X VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19620__A _19761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24878__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24461_ _25023_/CLK _24461_/D HRESETn VGND VGND VPWR VPWR _15032_/A sky130_fd_sc_hd__dfrtp_4
X_21673_ _21673_/A _20028_/Y VGND VGND VPWR VPWR _21674_/C sky130_fd_sc_hd__or2_4
XANTENNA__24807__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23412_ _23565_/CLK _23412_/D VGND VGND VPWR VPWR _20381_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_240_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20624_ _20624_/A _17413_/A VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__and2_4
X_24392_ _24378_/CLK _24392_/D HRESETn VGND VGND VPWR VPWR _17041_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23343_ _16550_/A _22485_/X _22852_/X _23342_/X VGND VGND VPWR VPWR _23344_/C sky130_fd_sc_hd__a211o_4
X_20555_ _20552_/A _20555_/B VGND VGND VPWR VPWR _20557_/B sky130_fd_sc_hd__nand2_4
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20359__A1_N _21991_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23274_ _24614_/Q _23274_/B VGND VGND VPWR VPWR _23274_/X sky130_fd_sc_hd__or2_4
X_20486_ _20486_/A VGND VGND VPWR VPWR _20486_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25013_ _25011_/CLK _15297_/X HRESETn VGND VGND VPWR VPWR _25013_/Q sky130_fd_sc_hd__dfrtp_4
X_22225_ _22209_/A _22223_/X _22224_/X VGND VGND VPWR VPWR _22229_/B sky130_fd_sc_hd__and3_4
XANTENNA__20799__A1 _15588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22156_ _21300_/Y VGND VGND VPWR VPWR _22157_/C sky130_fd_sc_hd__buf_2
XANTENNA__21460__A2 _21456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_219_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21107_ _21106_/X VGND VGND VPWR VPWR _21107_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22087_ _22387_/A _22087_/B _22087_/C VGND VGND VPWR VPWR _22087_/X sky130_fd_sc_hd__and3_4
XFILLER_247_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21038_ _22947_/A VGND VGND VPWR VPWR _22541_/A sky130_fd_sc_hd__buf_2
XANTENNA__18613__B1 _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22221__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13860_ _25258_/Q _13871_/A _13872_/A VGND VGND VPWR VPWR _13867_/A sky130_fd_sc_hd__or3_4
XFILLER_207_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12811_ _12858_/B VGND VGND VPWR VPWR _12912_/B sky130_fd_sc_hd__buf_2
XFILLER_16_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13791_ _21222_/B VGND VGND VPWR VPWR _13792_/A sky130_fd_sc_hd__buf_2
X_22989_ _24638_/Q _23165_/B VGND VGND VPWR VPWR _22989_/X sky130_fd_sc_hd__or2_4
XFILLER_231_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15530_ _11739_/B VGND VGND VPWR VPWR _15530_/Y sky130_fd_sc_hd__inv_2
X_12742_ _12742_/A _12738_/B VGND VGND VPWR VPWR _12742_/Y sky130_fd_sc_hd__nand2_4
X_24728_ _24732_/CLK _24728_/D HRESETn VGND VGND VPWR VPWR _16065_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_190_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _23946_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_187_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12673_ _12730_/A VGND VGND VPWR VPWR _12680_/A sky130_fd_sc_hd__buf_2
X_15461_ _15443_/A VGND VGND VPWR VPWR _15461_/X sky130_fd_sc_hd__buf_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _24169_/CLK _24659_/D HRESETn VGND VGND VPWR VPWR _22312_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_203_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24548__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17200_/A _17200_/B _17196_/X _17200_/D VGND VGND VPWR VPWR _17211_/C sky130_fd_sc_hd__or4_4
Xclkbuf_8_47_0_HCLK clkbuf_8_46_0_HCLK/A VGND VGND VPWR VPWR _23400_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14412_/A VGND VGND VPWR VPWR _14412_/X sky130_fd_sc_hd__buf_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18051_/A _18176_/X _18180_/C VGND VGND VPWR VPWR _18188_/B sky130_fd_sc_hd__or3_4
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _15142_/Y _15390_/A VGND VGND VPWR VPWR _15392_/X sky130_fd_sc_hd__or2_4
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17045_/A _17130_/Y VGND VGND VPWR VPWR _17131_/X sky130_fd_sc_hd__or2_4
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _25172_/Q _14342_/X _14334_/X VGND VGND VPWR VPWR _14343_/X sky130_fd_sc_hd__a21o_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14274_ _14272_/Y _14268_/X _13849_/X _14273_/X VGND VGND VPWR VPWR _14274_/X sky130_fd_sc_hd__a2bb2o_4
X_17062_ _17062_/A _17062_/B VGND VGND VPWR VPWR _17062_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13225_ _13315_/A _13225_/B _13224_/X VGND VGND VPWR VPWR _13225_/X sky130_fd_sc_hd__or3_4
X_16013_ _16010_/Y _16006_/X _15948_/X _16012_/X VGND VGND VPWR VPWR _16013_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13156_ _13155_/X VGND VGND VPWR VPWR _13178_/A sky130_fd_sc_hd__buf_2
XANTENNA__18852__B1 _16522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _12107_/A VGND VGND VPWR VPWR _12107_/X sky130_fd_sc_hd__buf_2
XFILLER_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13087_ _13087_/A VGND VGND VPWR VPWR _13087_/Y sky130_fd_sc_hd__inv_2
X_17964_ _17945_/A _17962_/X _17963_/X VGND VGND VPWR VPWR _17964_/X sky130_fd_sc_hd__and3_4
XFILLER_97_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19703_ _13288_/B VGND VGND VPWR VPWR _19703_/Y sky130_fd_sc_hd__inv_2
X_12038_ _12050_/A VGND VGND VPWR VPWR _12038_/X sky130_fd_sc_hd__buf_2
X_16915_ _22883_/A _24281_/Q _16130_/Y _16914_/Y VGND VGND VPWR VPWR _16922_/A sky130_fd_sc_hd__o22a_4
X_17895_ _21066_/A _17895_/B VGND VGND VPWR VPWR _17895_/X sky130_fd_sc_hd__or2_4
XFILLER_78_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19634_ _19631_/Y _19625_/X _19632_/X _19633_/X VGND VGND VPWR VPWR _23682_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16846_ _16853_/A VGND VGND VPWR VPWR _16846_/X sky130_fd_sc_hd__buf_2
XFILLER_226_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19565_ _19565_/A VGND VGND VPWR VPWR _19565_/X sky130_fd_sc_hd__buf_2
XFILLER_225_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16777_ _16776_/Y _16773_/X _15759_/X _16773_/X VGND VGND VPWR VPWR _24463_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13989_ _14027_/B VGND VGND VPWR VPWR _14028_/D sky130_fd_sc_hd__inv_2
XFILLER_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18516_ _18516_/A _18516_/B VGND VGND VPWR VPWR _18517_/B sky130_fd_sc_hd__or2_4
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15728_ _12555_/Y _15727_/X _11758_/X _15727_/X VGND VGND VPWR VPWR _15728_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19496_ _19483_/Y VGND VGND VPWR VPWR _19496_/X sky130_fd_sc_hd__buf_2
XANTENNA__24971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18447_ _24183_/Q VGND VGND VPWR VPWR _18531_/A sky130_fd_sc_hd__inv_2
X_15659_ _15651_/X _15659_/B VGND VGND VPWR VPWR _15659_/X sky130_fd_sc_hd__or2_4
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24900__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21074__A1_N _21747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18378_ _18377_/X VGND VGND VPWR VPWR _18379_/A sky130_fd_sc_hd__inv_2
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23112__D _23111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17329_ _17262_/Y _17326_/D VGND VGND VPWR VPWR _17330_/B sky130_fd_sc_hd__or2_4
XFILLER_193_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17895__A _21066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17343__B1 _17288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20340_ _20340_/A VGND VGND VPWR VPWR _20340_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18503__B _18710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21210__A _21210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20271_ _20269_/Y _20270_/X _20249_/X _20270_/X VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19096__B1 _18999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22010_ _22007_/Y _22008_/X _21996_/X _22009_/X VGND VGND VPWR VPWR _23358_/B sky130_fd_sc_hd__a211o_4
XFILLER_89_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23137__A _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23961_ _25223_/CLK _20606_/Y HRESETn VGND VGND VPWR VPWR _23961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22912_ _22487_/A _22911_/X VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__and2_4
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23892_ _23885_/CLK _23892_/D VGND VGND VPWR VPWR _23892_/Q sky130_fd_sc_hd__dfxtp_4
X_22843_ _20911_/C _22842_/X _20772_/C _22298_/A VGND VGND VPWR VPWR _22843_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22695__B _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22774_ _22757_/Y _22762_/Y _22770_/Y _21455_/X _22773_/X VGND VGND VPWR VPWR _22774_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_200_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24192_/CLK sky130_fd_sc_hd__clkbuf_1
X_21725_ _21293_/X _21711_/X _21714_/X _21721_/X _21724_/X VGND VGND VPWR VPWR _21841_/A
+ sky130_fd_sc_hd__o41a_4
X_24513_ _24073_/CLK _24513_/D HRESETn VGND VGND VPWR VPWR _24513_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25493_ _24196_/CLK _12054_/X HRESETn VGND VGND VPWR VPWR _25493_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24641__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11911__A RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_6_0_HCLK clkbuf_8_6_0_HCLK/A VGND VGND VPWR VPWR _23553_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14396__B1 _13846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21656_ _21972_/B VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__buf_2
X_24444_ _24476_/CLK _16819_/X HRESETn VGND VGND VPWR VPWR _24444_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21104__B _21104_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12946__A1 _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20607_ _14414_/Y _18893_/A _18876_/A _18890_/A VGND VGND VPWR VPWR _20608_/B sky130_fd_sc_hd__o22a_4
XFILLER_138_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24375_ _24639_/CLK _24375_/D HRESETn VGND VGND VPWR VPWR _24375_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21587_ _21565_/Y _21573_/X _21576_/X _21586_/Y VGND VGND VPWR VPWR _21610_/B sky130_fd_sc_hd__a211o_4
X_23326_ _21530_/X _23325_/X _21532_/X _15999_/A _21538_/X VGND VGND VPWR VPWR _23327_/A
+ sky130_fd_sc_hd__a32o_4
X_20538_ _24086_/Q _20543_/B _20526_/X VGND VGND VPWR VPWR _20538_/X sky130_fd_sc_hd__a21o_4
XFILLER_181_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14699__B2 _14761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23257_ _23188_/X _23254_/X _23256_/X VGND VGND VPWR VPWR _23258_/D sky130_fd_sc_hd__and3_4
X_20469_ _20469_/A _20469_/B VGND VGND VPWR VPWR _20469_/X sky130_fd_sc_hd__or2_4
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21969__B1 _21968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13010_ _13021_/A _13026_/C _13024_/A _13021_/D VGND VGND VPWR VPWR _13010_/X sky130_fd_sc_hd__or4_4
X_22208_ _21259_/A _20062_/Y VGND VGND VPWR VPWR _22209_/C sky130_fd_sc_hd__or2_4
XFILLER_165_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23188_ _22171_/A VGND VGND VPWR VPWR _23188_/X sky130_fd_sc_hd__buf_2
XFILLER_79_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15648__B1 _15489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22139_ _22139_/A _21719_/B VGND VGND VPWR VPWR _22139_/X sky130_fd_sc_hd__or2_4
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14961_ _15250_/A VGND VGND VPWR VPWR _14962_/A sky130_fd_sc_hd__inv_2
XFILLER_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16700_ _16699_/Y _16697_/X _15759_/X _16697_/X VGND VGND VPWR VPWR _16700_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13912_ _13915_/A VGND VGND VPWR VPWR _13955_/A sky130_fd_sc_hd__buf_2
X_17680_ _17585_/C _17683_/B _17600_/X VGND VGND VPWR VPWR _17680_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14892_ _14891_/X VGND VGND VPWR VPWR _25046_/D sky130_fd_sc_hd__inv_2
XFILLER_236_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14388__B _14388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16631_ _16631_/A VGND VGND VPWR VPWR _21167_/A sky130_fd_sc_hd__inv_2
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13843_ _13584_/Y _13838_/X _11838_/X _13842_/X VGND VGND VPWR VPWR _25268_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24729__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15820__B1 _11790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19350_ _18012_/B VGND VGND VPWR VPWR _19350_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16562_ _16562_/A VGND VGND VPWR VPWR _16562_/Y sky130_fd_sc_hd__inv_2
X_13774_ _13757_/C VGND VGND VPWR VPWR _13774_/X sky130_fd_sc_hd__buf_2
XFILLER_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18301_ _18301_/A _18301_/B VGND VGND VPWR VPWR _18301_/X sky130_fd_sc_hd__and2_4
X_15513_ _15503_/A VGND VGND VPWR VPWR _15513_/X sky130_fd_sc_hd__buf_2
XFILLER_31_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12725_ _12725_/A _12715_/X VGND VGND VPWR VPWR _12726_/C sky130_fd_sc_hd__nand2_4
X_19281_ _19280_/Y VGND VGND VPWR VPWR _19281_/X sky130_fd_sc_hd__buf_2
X_16493_ _16492_/Y _16488_/X _16407_/X _16488_/X VGND VGND VPWR VPWR _24574_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18232_ _18200_/A _19230_/A VGND VGND VPWR VPWR _18233_/C sky130_fd_sc_hd__or2_4
XFILLER_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11821__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15444_ _15444_/A _15447_/A VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__or2_4
XFILLER_31_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22449__A1 _12778_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _12630_/B _12647_/D _12630_/A VGND VGND VPWR VPWR _12656_/X sky130_fd_sc_hd__o21a_4
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22449__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ _18131_/A _18163_/B _18163_/C VGND VGND VPWR VPWR _18163_/X sky130_fd_sc_hd__or3_4
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _12587_/A _12582_/X _12584_/X _12586_/X VGND VGND VPWR VPWR _12608_/B sky130_fd_sc_hd__or4_4
X_15375_ _15306_/B _15381_/B VGND VGND VPWR VPWR _15376_/B sky130_fd_sc_hd__or2_4
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _17042_/B _17120_/B VGND VGND VPWR VPWR _17115_/B sky130_fd_sc_hd__or2_4
XANTENNA__14139__B1 _14137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _25179_/Q _14308_/Y _25178_/Q _14316_/A VGND VGND VPWR VPWR _14326_/X sky130_fd_sc_hd__o22a_4
X_18094_ _18200_/A _23897_/Q VGND VGND VPWR VPWR _18095_/C sky130_fd_sc_hd__or2_4
XFILLER_209_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17045_ _17045_/A VGND VGND VPWR VPWR _17132_/A sky130_fd_sc_hd__inv_2
XANTENNA__13748__A _13748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14257_ _13949_/Y _13958_/X _13969_/Y _14257_/D VGND VGND VPWR VPWR _14257_/X sky130_fd_sc_hd__or4_4
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13208_ _13208_/A VGND VGND VPWR VPWR _13209_/A sky130_fd_sc_hd__inv_2
X_14188_ _14186_/Y _14119_/X _14145_/X _14187_/Y VGND VGND VPWR VPWR _14188_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15639__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15963__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13139_ _13139_/A _13138_/X VGND VGND VPWR VPWR _13139_/X sky130_fd_sc_hd__or2_4
XFILLER_124_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19435__A _17963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18996_ _18996_/A VGND VGND VPWR VPWR _18996_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17947_ _17943_/A _19141_/A VGND VGND VPWR VPWR _17947_/X sky130_fd_sc_hd__or2_4
XFILLER_39_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19250__B1 _19226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17878_ _16920_/Y _17877_/X _16964_/X VGND VGND VPWR VPWR _17878_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16064__B1 _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16829_ _14936_/Y _16825_/X HWDATA[19] _16828_/X VGND VGND VPWR VPWR _16829_/X sky130_fd_sc_hd__a2bb2o_4
X_19617_ _19617_/A VGND VGND VPWR VPWR _21976_/B sky130_fd_sc_hd__inv_2
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22137__B1 _22105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19548_ _19548_/A _14201_/A VGND VGND VPWR VPWR _21217_/A sky130_fd_sc_hd__or2_4
XANTENNA__22688__A1 _16244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19479_ _19479_/A VGND VGND VPWR VPWR _22357_/B sky130_fd_sc_hd__inv_2
X_21510_ _21278_/X VGND VGND VPWR VPWR _22400_/A sky130_fd_sc_hd__buf_2
X_22490_ _22490_/A _22985_/B VGND VGND VPWR VPWR _22490_/X sky130_fd_sc_hd__or2_4
XANTENNA__24052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_30_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24386_/CLK sky130_fd_sc_hd__clkbuf_1
X_21441_ _21440_/X VGND VGND VPWR VPWR _21711_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_93_0_HCLK clkbuf_7_46_0_HCLK/X VGND VGND VPWR VPWR _25425_/CLK sky130_fd_sc_hd__clkbuf_1
X_24160_ _24160_/CLK _24160_/D HRESETn VGND VGND VPWR VPWR _24160_/Q sky130_fd_sc_hd__dfrtp_4
X_21372_ _25250_/Q VGND VGND VPWR VPWR _21372_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14761__B _14753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23111_ _23106_/Y _23110_/Y _22868_/X VGND VGND VPWR VPWR _23111_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15878__B1 _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20323_ _20323_/A VGND VGND VPWR VPWR _20323_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24091_ _24966_/CLK _24091_/D HRESETn VGND VGND VPWR VPWR _20487_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__19069__B1 _18975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23042_ _23106_/A _23041_/X VGND VGND VPWR VPWR _23042_/Y sky130_fd_sc_hd__nor2_4
X_20254_ _20253_/Y _20248_/X _19761_/X _20234_/Y VGND VGND VPWR VPWR _23461_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20185_ _20183_/Y _20184_/X _20119_/X _20184_/X VGND VGND VPWR VPWR _23487_/D sky130_fd_sc_hd__a2bb2o_4
X_24993_ _24975_/CLK _24993_/D HRESETn VGND VGND VPWR VPWR _24993_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23944_ _24095_/CLK _23944_/D HRESETn VGND VGND VPWR VPWR _20998_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24893__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23875_ _23871_/CLK _19080_/X VGND VGND VPWR VPWR _13213_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_217_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24822__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22826_ _22944_/A VGND VGND VPWR VPWR _23025_/A sky130_fd_sc_hd__buf_2
XANTENNA__22679__A1 _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25545_ _24327_/CLK _25545_/D HRESETn VGND VGND VPWR VPWR _25545_/Q sky130_fd_sc_hd__dfrtp_4
X_22757_ _21060_/A _22757_/B VGND VGND VPWR VPWR _22757_/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12510_ _12273_/X _12508_/X _12509_/Y VGND VGND VPWR VPWR _25441_/D sky130_fd_sc_hd__o21a_4
X_13490_ _13490_/A VGND VGND VPWR VPWR _13490_/Y sky130_fd_sc_hd__inv_2
X_21708_ _21557_/X _21610_/X _21708_/C _21707_/X VGND VGND VPWR VPWR HRDATA[2] sky130_fd_sc_hd__or4_4
X_22688_ _16244_/Y _22462_/X _16430_/Y _22459_/X VGND VGND VPWR VPWR _22689_/B sky130_fd_sc_hd__o22a_4
X_25476_ _24196_/CLK _12129_/X HRESETn VGND VGND VPWR VPWR _25476_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12919__A1 _12834_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12441_ _12295_/X _12449_/D VGND VGND VPWR VPWR _12442_/B sky130_fd_sc_hd__or2_4
X_21639_ _22388_/A _19873_/Y VGND VGND VPWR VPWR _21639_/X sky130_fd_sc_hd__or2_4
X_24427_ _24425_/CLK _24427_/D HRESETn VGND VGND VPWR VPWR _14925_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_139_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13041__B1 _13040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17307__B1 _17288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _12372_/A VGND VGND VPWR VPWR _13004_/B sky130_fd_sc_hd__inv_2
X_15160_ _25003_/Q _15158_/Y _15362_/A _24605_/Q VGND VGND VPWR VPWR _15161_/D sky130_fd_sc_hd__a2bb2o_4
X_24358_ _24346_/CLK _17352_/Y HRESETn VGND VGND VPWR VPWR _17258_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_1_0_HCLK clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14111_ _14111_/A _14111_/B _25226_/Q VGND VGND VPWR VPWR _14112_/B sky130_fd_sc_hd__or3_4
X_15091_ _15091_/A _15085_/X _15091_/C _15091_/D VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__or4_4
X_23309_ _23309_/A _22849_/X VGND VGND VPWR VPWR _23309_/X sky130_fd_sc_hd__or2_4
X_24289_ _24272_/CLK _17801_/Y HRESETn VGND VGND VPWR VPWR _24289_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12472__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14042_ _25247_/Q _14042_/B VGND VGND VPWR VPWR _14042_/X sky130_fd_sc_hd__or2_4
XFILLER_107_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18850_ _18846_/X _18850_/B _18850_/C _18849_/X VGND VGND VPWR VPWR _18850_/X sky130_fd_sc_hd__or4_4
XFILLER_122_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17801_ _17801_/A VGND VGND VPWR VPWR _17801_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18781_ _18780_/X VGND VGND VPWR VPWR _18782_/B sky130_fd_sc_hd__inv_2
X_15993_ _11861_/A VGND VGND VPWR VPWR _15993_/X sky130_fd_sc_hd__buf_2
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19298__A2_N _19293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17732_ _17732_/A VGND VGND VPWR VPWR _17732_/X sky130_fd_sc_hd__buf_2
XFILLER_248_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14944_ _15270_/A _24428_/Q _15271_/A _14943_/Y VGND VGND VPWR VPWR _14948_/C sky130_fd_sc_hd__o22a_4
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17663_ _17663_/A _17589_/X VGND VGND VPWR VPWR _17664_/B sky130_fd_sc_hd__or2_4
XFILLER_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14875_ _14875_/A VGND VGND VPWR VPWR _14875_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24563__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21590__A1 _14946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19402_ _19131_/A VGND VGND VPWR VPWR _19402_/X sky130_fd_sc_hd__buf_2
XFILLER_223_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _16612_/Y _16610_/X _16613_/X _16610_/X VGND VGND VPWR VPWR _16614_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13826_ _21280_/A VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__buf_2
XANTENNA__15550__A2_N _15547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17594_ _17663_/A _17525_/Y _17569_/X _17594_/D VGND VGND VPWR VPWR _17595_/B sky130_fd_sc_hd__or4_4
XFILLER_235_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19333_ _23785_/Q VGND VGND VPWR VPWR _19333_/Y sky130_fd_sc_hd__inv_2
X_16545_ _16544_/Y _16540_/X _16451_/X _16540_/X VGND VGND VPWR VPWR _16545_/X sky130_fd_sc_hd__a2bb2o_4
X_13757_ _13757_/A _13772_/A _13757_/C _25284_/Q VGND VGND VPWR VPWR _13757_/X sky130_fd_sc_hd__and4_4
X_12708_ _12574_/Y _12702_/X _12705_/B _12662_/X VGND VGND VPWR VPWR _12708_/X sky130_fd_sc_hd__a211o_4
X_19264_ _19258_/Y VGND VGND VPWR VPWR _19264_/X sky130_fd_sc_hd__buf_2
X_16476_ _16495_/A VGND VGND VPWR VPWR _16476_/X sky130_fd_sc_hd__buf_2
XFILLER_188_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13688_ _13703_/B VGND VGND VPWR VPWR _13688_/Y sky130_fd_sc_hd__inv_2
X_18215_ _14656_/A _18213_/X _18215_/C VGND VGND VPWR VPWR _18215_/X sky130_fd_sc_hd__and3_4
X_15427_ _15425_/Y _15426_/X _15427_/C VGND VGND VPWR VPWR _15427_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_34_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12639_ _12631_/X _12647_/D _12601_/Y VGND VGND VPWR VPWR _12640_/C sky130_fd_sc_hd__o21a_4
X_19195_ _19195_/A VGND VGND VPWR VPWR _19195_/Y sky130_fd_sc_hd__inv_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18146_ _17987_/A _20247_/A VGND VGND VPWR VPWR _18146_/X sky130_fd_sc_hd__or2_4
X_15358_ _15358_/A VGND VGND VPWR VPWR _25003_/D sky130_fd_sc_hd__inv_2
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14309_ _14309_/A _14308_/Y VGND VGND VPWR VPWR _14310_/C sky130_fd_sc_hd__or2_4
XANTENNA__25351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18077_ _17987_/A _23465_/Q VGND VGND VPWR VPWR _18077_/X sky130_fd_sc_hd__or2_4
X_15289_ _14990_/X _15291_/B _15288_/Y VGND VGND VPWR VPWR _15289_/X sky130_fd_sc_hd__o21a_4
X_17028_ _17355_/B VGND VGND VPWR VPWR _17345_/A sky130_fd_sc_hd__buf_2
XANTENNA__19471__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18979_ _18979_/A VGND VGND VPWR VPWR _18979_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19223__B1 _19131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21990_ _18372_/A _20360_/Y _18357_/A _21991_/B VGND VGND VPWR VPWR _21990_/X sky130_fd_sc_hd__o22a_4
XFILLER_227_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16037__B1 _15967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20941_ _20944_/B _13674_/X _20940_/Y VGND VGND VPWR VPWR _20941_/Y sky130_fd_sc_hd__a21oi_4
XPHY_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12133__A1_N _12132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17413__A _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20872_ _16708_/Y _20854_/X _20863_/X _20871_/Y VGND VGND VPWR VPWR _20872_/X sky130_fd_sc_hd__o22a_4
X_23660_ _23916_/CLK _19700_/X VGND VGND VPWR VPWR _13162_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22611_ _22289_/A _22610_/X _21314_/X _24732_/Q _21317_/X VGND VGND VPWR VPWR _22611_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _23590_/CLK _23591_/D VGND VGND VPWR VPWR _23591_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22542_ _22542_/A VGND VGND VPWR VPWR _22542_/X sky130_fd_sc_hd__buf_2
X_25330_ _25494_/CLK _25330_/D HRESETn VGND VGND VPWR VPWR _13474_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22473_ _21606_/X VGND VGND VPWR VPWR _22476_/A sky130_fd_sc_hd__buf_2
X_25261_ _25276_/CLK _25261_/D HRESETn VGND VGND VPWR VPWR _25261_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15868__A _23053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21424_ _21423_/X VGND VGND VPWR VPWR _21425_/D sky130_fd_sc_hd__inv_2
X_24212_ _23459_/CLK _24212_/D HRESETn VGND VGND VPWR VPWR _17478_/B sky130_fd_sc_hd__dfrtp_4
X_25192_ _25253_/CLK _25192_/D HRESETn VGND VGND VPWR VPWR _25192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24143_ _24145_/CLK _18786_/Y HRESETn VGND VGND VPWR VPWR _18693_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13388__A _13420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21355_ _14186_/Y _22334_/B _23938_/Q _21369_/B VGND VGND VPWR VPWR _21361_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20306_ _22268_/B _20303_/X _19993_/X _20303_/X VGND VGND VPWR VPWR _23442_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24074_ _24503_/CLK _24074_/D HRESETn VGND VGND VPWR VPWR _24074_/Q sky130_fd_sc_hd__dfrtp_4
X_21286_ _18277_/X _21284_/X _21180_/X _21285_/Y VGND VGND VPWR VPWR _21286_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23025_ _23025_/A _23025_/B _23025_/C VGND VGND VPWR VPWR _23025_/X sky130_fd_sc_hd__and3_4
XFILLER_116_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20237_ _17987_/B VGND VGND VPWR VPWR _20237_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19462__B1 _19439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20168_ _21273_/B _20163_/X _20146_/X _20150_/Y VGND VGND VPWR VPWR _20168_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_218_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12990_ _21056_/A _12875_/X _12989_/Y VGND VGND VPWR VPWR _12990_/X sky130_fd_sc_hd__o21a_4
X_20099_ _20099_/A VGND VGND VPWR VPWR _20099_/Y sky130_fd_sc_hd__inv_2
X_24976_ _24979_/CLK _15452_/X HRESETn VGND VGND VPWR VPWR _13934_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11941_ _19996_/A VGND VGND VPWR VPWR _19632_/A sky130_fd_sc_hd__buf_2
X_23927_ _23926_/CLK _23927_/D VGND VGND VPWR VPWR _23927_/Q sky130_fd_sc_hd__dfxtp_4
X_14660_ _18013_/A VGND VGND VPWR VPWR _17944_/A sky130_fd_sc_hd__buf_2
XFILLER_232_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11872_ _11869_/Y _11750_/X _11871_/X _11750_/X VGND VGND VPWR VPWR _25526_/D sky130_fd_sc_hd__a2bb2o_4
X_23858_ _23871_/CLK _19127_/X VGND VGND VPWR VPWR _13272_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_221_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13611_ _13611_/A VGND VGND VPWR VPWR _19346_/B sky130_fd_sc_hd__buf_2
X_22809_ _20772_/A _22298_/X _20906_/Y _22808_/X VGND VGND VPWR VPWR _22809_/X sky130_fd_sc_hd__o22a_4
XFILLER_232_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14591_ _14586_/C _14588_/X VGND VGND VPWR VPWR _14591_/X sky130_fd_sc_hd__or2_4
XFILLER_198_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23789_ _23794_/CLK _23789_/D VGND VGND VPWR VPWR _13460_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16330_ _16329_/Y _16325_/X _15972_/X _16325_/X VGND VGND VPWR VPWR _16330_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13542_ _13484_/C _13484_/D _13542_/C _12109_/A VGND VGND VPWR VPWR _13543_/A sky130_fd_sc_hd__or4_4
X_25528_ _25528_/CLK _25528_/D HRESETn VGND VGND VPWR VPWR _25528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16200__B1 _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16261_ _22312_/A VGND VGND VPWR VPWR _16261_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13473_ _13207_/A _13472_/X _25331_/Q _13267_/A VGND VGND VPWR VPWR _13473_/X sky130_fd_sc_hd__o22a_4
X_25459_ _25456_/CLK _25459_/D HRESETn VGND VGND VPWR VPWR _12293_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18000_ _18008_/A VGND VGND VPWR VPWR _18158_/A sky130_fd_sc_hd__buf_2
X_15212_ _14964_/A _15215_/B VGND VGND VPWR VPWR _15213_/C sky130_fd_sc_hd__or2_4
X_12424_ _12424_/A _12424_/B VGND VGND VPWR VPWR _12425_/B sky130_fd_sc_hd__or2_4
XANTENNA__25109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16192_ _16192_/A VGND VGND VPWR VPWR _22462_/A sky130_fd_sc_hd__buf_2
XFILLER_154_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15143_ _15142_/Y _16430_/A _15142_/Y _16430_/A VGND VGND VPWR VPWR _15143_/X sky130_fd_sc_hd__a2bb2o_4
X_12355_ _13003_/A _12353_/Y _12351_/A _12354_/Y VGND VGND VPWR VPWR _12355_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _12428_/A _12425_/A VGND VGND VPWR VPWR _12298_/C sky130_fd_sc_hd__or2_4
X_15074_ _15074_/A VGND VGND VPWR VPWR _15075_/C sky130_fd_sc_hd__inv_2
X_19951_ _19958_/A VGND VGND VPWR VPWR _19951_/X sky130_fd_sc_hd__buf_2
XANTENNA__15857__A3 _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14025_ _13994_/A _13994_/B VGND VGND VPWR VPWR _14025_/Y sky130_fd_sc_hd__nand2_4
X_18902_ _14388_/B _17450_/B VGND VGND VPWR VPWR _18902_/Y sky130_fd_sc_hd__nor2_4
X_19882_ _19882_/A VGND VGND VPWR VPWR _19895_/A sky130_fd_sc_hd__inv_2
XANTENNA__16402__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16267__B1 _16073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18833_ _16546_/Y _24132_/Q _24557_/Q _18809_/A VGND VGND VPWR VPWR _18833_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24744__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18764_ _18764_/A _18764_/B VGND VGND VPWR VPWR _18769_/B sky130_fd_sc_hd__or2_4
X_15976_ _15974_/X _15943_/X HWDATA[16] _22778_/A _15975_/X VGND VGND VPWR VPWR _24769_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_209_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17715_ _21212_/A VGND VGND VPWR VPWR _17716_/A sky130_fd_sc_hd__buf_2
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14927_ _14927_/A VGND VGND VPWR VPWR _15203_/A sky130_fd_sc_hd__inv_2
X_18695_ _24145_/Q VGND VGND VPWR VPWR _18772_/A sky130_fd_sc_hd__inv_2
XFILLER_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17646_ _17531_/Y _17578_/B _17646_/C _17646_/D VGND VGND VPWR VPWR _17652_/B sky130_fd_sc_hd__or4_4
XFILLER_224_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14858_ _25054_/Q _14810_/B _25054_/Q _14810_/B VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13809_ _14412_/A VGND VGND VPWR VPWR _13809_/X sky130_fd_sc_hd__buf_2
X_17577_ _17516_/Y _17646_/C _17577_/C _17644_/A VGND VGND VPWR VPWR _17577_/X sky130_fd_sc_hd__or4_4
X_14789_ _14789_/A VGND VGND VPWR VPWR _14789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17519__B1 _11837_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22512__B1 _21591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19316_ _19301_/Y VGND VGND VPWR VPWR _19316_/X sky130_fd_sc_hd__buf_2
X_16528_ _16527_/Y _16525_/X _16157_/X _16525_/X VGND VGND VPWR VPWR _16528_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19247_ _19245_/Y _19241_/X _19246_/X _19241_/X VGND VGND VPWR VPWR _19247_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16459_ _23009_/A VGND VGND VPWR VPWR _16460_/A sky130_fd_sc_hd__buf_2
XANTENNA__17179__A1_N _24623_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18064__A _18098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19178_ _18133_/B VGND VGND VPWR VPWR _19178_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18999__A _19139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18129_ _18129_/A _23896_/Q VGND VGND VPWR VPWR _18130_/C sky130_fd_sc_hd__or2_4
XFILLER_117_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_104_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24639_/CLK sky130_fd_sc_hd__clkbuf_1
X_21140_ _21140_/A _17448_/C _14415_/A _13822_/B VGND VGND VPWR VPWR _21353_/A sky130_fd_sc_hd__or4_4
XFILLER_105_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_167_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23522_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21071_ _21071_/A _15667_/A VGND VGND VPWR VPWR _21071_/X sky130_fd_sc_hd__and2_4
XANTENNA__16258__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20022_ _20016_/Y VGND VGND VPWR VPWR _20022_/X sky130_fd_sc_hd__buf_2
XFILLER_247_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22968__B _22968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24830_ _24849_/CLK _24830_/D HRESETn VGND VGND VPWR VPWR _24830_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24761_ _24759_/CLK _24761_/D HRESETn VGND VGND VPWR VPWR _12213_/A sky130_fd_sc_hd__dfrtp_4
X_21973_ _18268_/X _21971_/X _21972_/X _13795_/Y _21654_/X VGND VGND VPWR VPWR _21974_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_66_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13492__B1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21554__B2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23712_ _23407_/CLK _19539_/X VGND VGND VPWR VPWR _19538_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _20923_/Y _20924_/B VGND VGND VPWR VPWR _20924_/X sky130_fd_sc_hd__and2_4
XFILLER_242_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24692_ _24689_/CLK _24692_/D HRESETn VGND VGND VPWR VPWR _22201_/A sky130_fd_sc_hd__dfrtp_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _13666_/A VGND VGND VPWR VPWR _20855_/Y sky130_fd_sc_hd__inv_2
X_23643_ _23644_/CLK _23643_/D VGND VGND VPWR VPWR _13258_/B sky130_fd_sc_hd__dfxtp_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _20790_/B _20779_/X _20785_/X VGND VGND VPWR VPWR _20786_/Y sky130_fd_sc_hd__a21oi_4
X_23574_ _23597_/CLK _19941_/X VGND VGND VPWR VPWR _19940_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25313_ _25188_/CLK _13525_/X HRESETn VGND VGND VPWR VPWR _13523_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22525_ _22525_/A _22468_/X VGND VGND VPWR VPWR _22525_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14933__C _14929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25244_ _25105_/CLK _14083_/X HRESETn VGND VGND VPWR VPWR _25244_/Q sky130_fd_sc_hd__dfrtp_4
X_22456_ _17364_/B _22442_/A _25446_/Q _22487_/A VGND VGND VPWR VPWR _22458_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21407_ _14688_/X _21407_/B VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__or2_4
X_22387_ _22387_/A _22387_/B _22387_/C VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__and3_4
X_25175_ _23954_/CLK _25175_/D HRESETn VGND VGND VPWR VPWR _25175_/Q sky130_fd_sc_hd__dfrtp_4
X_12140_ _12140_/A _20982_/A VGND VGND VPWR VPWR _12140_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__23965__D sda_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21338_ _22171_/A _21338_/B _21338_/C VGND VGND VPWR VPWR _21338_/X sky130_fd_sc_hd__and3_4
X_24126_ _23946_/CLK _24126_/D HRESETn VGND VGND VPWR VPWR _24126_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_151_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12055_/Y _12070_/Y _11876_/X _12070_/Y VGND VGND VPWR VPWR _25492_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13846__A _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21269_ _21265_/X _21268_/X _21251_/X VGND VGND VPWR VPWR _21269_/X sky130_fd_sc_hd__o21a_4
X_24057_ _24493_/CLK _24057_/D HRESETn VGND VGND VPWR VPWR _24057_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23039__B _23036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16249__B1 _16248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23008_ _23008_/A _23007_/X VGND VGND VPWR VPWR _23008_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22878__B _22789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15830_ _15825_/X _15828_/X _15754_/X _24839_/Q _15826_/X VGND VGND VPWR VPWR _15830_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15761_ HWDATA[11] VGND VGND VPWR VPWR _15761_/X sky130_fd_sc_hd__buf_2
XFILLER_246_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12973_ _12984_/A _12969_/X _12972_/Y VGND VGND VPWR VPWR _25379_/D sky130_fd_sc_hd__and3_4
X_24959_ _23991_/CLK _15484_/X HRESETn VGND VGND VPWR VPWR _24959_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_206_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21545__A1 _15565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17500_ _17490_/Y _17491_/X _17492_/X _17499_/X VGND VGND VPWR VPWR _17500_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21545__B2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14712_ _14712_/A _14713_/A _14707_/X _14711_/X VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__or4_4
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11924_ _11886_/A _11923_/X _11921_/Y VGND VGND VPWR VPWR _25518_/D sky130_fd_sc_hd__o21a_4
X_18480_ _24167_/Q VGND VGND VPWR VPWR _18480_/Y sky130_fd_sc_hd__inv_2
X_15692_ _15691_/X VGND VGND VPWR VPWR _15692_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17431_ _17429_/Y _17426_/X _17430_/X _17426_/X VGND VGND VPWR VPWR _17431_/X sky130_fd_sc_hd__a2bb2o_4
X_14643_ _14626_/A VGND VGND VPWR VPWR _14643_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11855_ _11855_/A VGND VGND VPWR VPWR _14400_/A sky130_fd_sc_hd__buf_2
XFILLER_221_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17362_ _17362_/A _17360_/A VGND VGND VPWR VPWR _17362_/X sky130_fd_sc_hd__or2_4
X_14574_ _14607_/A _14574_/B VGND VGND VPWR VPWR _14574_/X sky130_fd_sc_hd__or2_4
XFILLER_82_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ _11759_/X VGND VGND VPWR VPWR _11786_/X sky130_fd_sc_hd__buf_2
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19101_ _22379_/B _19100_/X _16872_/X _19100_/X VGND VGND VPWR VPWR _23868_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ _16311_/Y _16305_/X _15957_/X _16312_/X VGND VGND VPWR VPWR _24641_/D sky130_fd_sc_hd__a2bb2o_4
X_13525_ _13536_/A _13521_/X _13524_/X _13521_/X VGND VGND VPWR VPWR _13525_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17293_ _17293_/A _17292_/Y VGND VGND VPWR VPWR _17295_/B sky130_fd_sc_hd__or2_4
XANTENNA__12925__A _12819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19032_ _19032_/A VGND VGND VPWR VPWR _19032_/X sky130_fd_sc_hd__buf_2
X_16244_ _16244_/A VGND VGND VPWR VPWR _16244_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15301__A _15388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13456_ _13456_/A _13448_/X _13456_/C VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__and3_4
XFILLER_174_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12407_ _12409_/B VGND VGND VPWR VPWR _12408_/B sky130_fd_sc_hd__inv_2
X_16175_ _21069_/A VGND VGND VPWR VPWR _16175_/Y sky130_fd_sc_hd__inv_2
X_13387_ _13387_/A _13385_/X _13387_/C VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__and3_4
XANTENNA__24996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ _24999_/Q VGND VGND VPWR VPWR _15376_/A sky130_fd_sc_hd__inv_2
X_12338_ _13023_/A _24854_/Q _13024_/A _12337_/Y VGND VGND VPWR VPWR _12348_/A sky130_fd_sc_hd__o22a_4
XFILLER_115_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15057_ _14895_/X _24462_/Q _25017_/Q _15036_/Y VGND VGND VPWR VPWR _15057_/X sky130_fd_sc_hd__a2bb2o_4
X_19934_ _19933_/Y _19931_/X _19800_/X _19931_/X VGND VGND VPWR VPWR _19934_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12269_ _25458_/Q VGND VGND VPWR VPWR _12269_/Y sky130_fd_sc_hd__inv_2
X_14008_ _25246_/Q VGND VGND VPWR VPWR _14008_/X sky130_fd_sc_hd__buf_2
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_17_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19865_ _22218_/B _19862_/X _19793_/X _19862_/X VGND VGND VPWR VPWR _19865_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18816_ _24136_/Q _18815_/Y VGND VGND VPWR VPWR _18816_/X sky130_fd_sc_hd__or2_4
XFILLER_96_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19796_ _16874_/X VGND VGND VPWR VPWR _19796_/X sky130_fd_sc_hd__buf_2
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15959_ _15938_/X _15943_/X HWDATA[23] _23049_/A _15941_/X VGND VGND VPWR VPWR _24776_/D
+ sky130_fd_sc_hd__a32o_4
X_18747_ _18714_/A _18744_/B _18746_/X VGND VGND VPWR VPWR _18748_/A sky130_fd_sc_hd__or3_4
XFILLER_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12277__B2 _24757_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18059__A _18059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22733__B1 _24839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18678_ _24161_/Q VGND VGND VPWR VPWR _18678_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17629_ _24319_/Q _17629_/B VGND VGND VPWR VPWR _17630_/C sky130_fd_sc_hd__or2_4
XANTENNA__17898__A _17710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20640_ _15476_/Y _20623_/X _20637_/X _20639_/X VGND VGND VPWR VPWR _20640_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14974__B1 _25023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11788__B1 _11787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20571_ _20571_/A _20570_/Y _20556_/X VGND VGND VPWR VPWR _20571_/X sky130_fd_sc_hd__and3_4
X_22310_ _23299_/A _22301_/Y _22305_/X _22150_/A _22309_/X VGND VGND VPWR VPWR _22310_/X
+ sky130_fd_sc_hd__o32a_4
X_23290_ _23290_/A _23322_/B VGND VGND VPWR VPWR _23290_/X sky130_fd_sc_hd__or2_4
XFILLER_192_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22241_ _13560_/Y _22595_/B _21180_/X VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__a21o_4
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19665__B1 _19612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12201__B2 _24779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16479__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22172_ _16263_/A _22316_/B VGND VGND VPWR VPWR _22172_/X sky130_fd_sc_hd__or2_4
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24666__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21123_ _21123_/A VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__buf_2
XFILLER_105_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22979__A _22956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21054_ _21589_/B VGND VGND VPWR VPWR _21882_/A sky130_fd_sc_hd__buf_2
XFILLER_87_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20005_ _23551_/Q VGND VGND VPWR VPWR _21688_/B sky130_fd_sc_hd__inv_2
XANTENNA__22972__B1 _12375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_HCLK clkbuf_3_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24813_ _24856_/CLK _24813_/D HRESETn VGND VGND VPWR VPWR _23054_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14497__A _14485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24744_ _24372_/CLK _16027_/X HRESETn VGND VGND VPWR VPWR _24744_/Q sky130_fd_sc_hd__dfrtp_4
X_21956_ _21476_/A _21956_/B VGND VGND VPWR VPWR _21957_/C sky130_fd_sc_hd__or2_4
XFILLER_243_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _24063_/Q _20907_/B VGND VGND VPWR VPWR _20907_/X sky130_fd_sc_hd__or2_4
XFILLER_43_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24675_ _24674_/CLK _16218_/X HRESETn VGND VGND VPWR VPWR _23076_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _24757_/Q _21043_/A _22684_/B _24829_/Q _15553_/X VGND VGND VPWR VPWR _21887_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23628_/CLK _23626_/D VGND VGND VPWR VPWR _19795_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20837_/X VGND VGND VPWR VPWR _20838_/Y sky130_fd_sc_hd__inv_2
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23557_ _23565_/CLK _23557_/D VGND VGND VPWR VPWR _19983_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_10_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20769_ _20772_/A _20763_/Y _20768_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__o21a_4
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13164_/Y VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__buf_2
XFILLER_128_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _12229_/X _22507_/X _17871_/A _21079_/A VGND VGND VPWR VPWR _22508_/X sky130_fd_sc_hd__a2bb2o_4
X_14290_ _14290_/A VGND VGND VPWR VPWR _20684_/A sky130_fd_sc_hd__buf_2
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _23488_/CLK _23488_/D VGND VGND VPWR VPWR _23488_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13182_/A VGND VGND VPWR VPWR _13241_/X sky130_fd_sc_hd__buf_2
X_25227_ _23395_/CLK _14147_/X HRESETn VGND VGND VPWR VPWR _14112_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22439_ _22897_/A VGND VGND VPWR VPWR _22543_/A sky130_fd_sc_hd__buf_2
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19528__A _19527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13172_ _13163_/X _13169_/X _13171_/X VGND VGND VPWR VPWR _13172_/X sky130_fd_sc_hd__o21a_4
X_25158_ _24012_/CLK _25158_/D HRESETn VGND VGND VPWR VPWR _20477_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_170_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12123_ _12123_/A VGND VGND VPWR VPWR _12123_/X sky130_fd_sc_hd__buf_2
X_24109_ _23647_/CLK _20977_/X HRESETn VGND VGND VPWR VPWR _24109_/Q sky130_fd_sc_hd__dfrtp_4
X_17980_ _17975_/X _17977_/X _17979_/X VGND VGND VPWR VPWR _17980_/X sky130_fd_sc_hd__and3_4
XFILLER_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19408__B1 _19341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25089_ _25276_/CLK _25089_/D HRESETn VGND VGND VPWR VPWR _13561_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_150_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _25494_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22889__A _22887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12911__C _12609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12054_ _24111_/Q _12036_/X _25493_/Q _12050_/X VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__o22a_4
X_16931_ _16924_/X _16926_/X _16928_/X _16931_/D VGND VGND VPWR VPWR _16931_/X sky130_fd_sc_hd__or4_4
XFILLER_151_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16862_ _14946_/Y _16857_/X _16861_/X _16857_/X VGND VGND VPWR VPWR _16862_/X sky130_fd_sc_hd__a2bb2o_4
X_19650_ _23676_/Q VGND VGND VPWR VPWR _19650_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18631__A1 _16615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22401__B _22319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15813_ _15790_/X _15804_/X _15732_/X _24851_/Q _15802_/X VGND VGND VPWR VPWR _15813_/X
+ sky130_fd_sc_hd__a32o_4
X_18601_ _18597_/B _18600_/X _18598_/C VGND VGND VPWR VPWR _18601_/X sky130_fd_sc_hd__and3_4
XFILLER_65_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19581_ _22041_/B _19575_/X _11948_/X _19580_/X VGND VGND VPWR VPWR _23698_/D sky130_fd_sc_hd__a2bb2o_4
X_16793_ _15036_/Y _16787_/X _16791_/X _16792_/X VGND VGND VPWR VPWR _24455_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18532_ _18534_/B VGND VGND VPWR VPWR _18533_/B sky130_fd_sc_hd__inv_2
X_15744_ _15726_/X VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__buf_2
X_12956_ _12851_/A _12956_/B VGND VGND VPWR VPWR _12957_/C sky130_fd_sc_hd__or2_4
XFILLER_233_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18395__B1 _24196_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22191__B2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11907_ _11900_/A _11906_/Y _11902_/A VGND VGND VPWR VPWR _11907_/X sky130_fd_sc_hd__o21a_4
X_18463_ _18445_/Y _18510_/A VGND VGND VPWR VPWR _18488_/C sky130_fd_sc_hd__or2_4
XFILLER_34_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15675_ _21574_/A VGND VGND VPWR VPWR _15676_/A sky130_fd_sc_hd__buf_2
XFILLER_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12887_ _12886_/X VGND VGND VPWR VPWR _12888_/B sky130_fd_sc_hd__inv_2
XFILLER_206_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17414_ _17396_/X _17410_/X _24344_/Q _21010_/A _17413_/X VGND VGND VPWR VPWR _24345_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14626_/A _14626_/B VGND VGND VPWR VPWR _14626_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__25124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11838_ HWDATA[8] VGND VGND VPWR VPWR _11838_/X sky130_fd_sc_hd__buf_2
X_18394_ _18393_/Y _18391_/X _24196_/Q _18391_/X VGND VGND VPWR VPWR _24197_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/A _17256_/X VGND VGND VPWR VPWR _17345_/X sky130_fd_sc_hd__or2_4
XANTENNA__21033__A _21032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A VGND VGND VPWR VPWR _14557_/Y sky130_fd_sc_hd__inv_2
X_11769_ _11759_/X VGND VGND VPWR VPWR _11769_/X sky130_fd_sc_hd__buf_2
XFILLER_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _12032_/Y _13507_/X _11834_/X _13507_/X VGND VGND VPWR VPWR _13508_/X sky130_fd_sc_hd__a2bb2o_4
X_17276_ _17355_/B _17240_/X VGND VGND VPWR VPWR _17276_/X sky130_fd_sc_hd__and2_4
X_14488_ _14487_/Y _14485_/X _14423_/X _14485_/X VGND VGND VPWR VPWR _25125_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19015_ _23897_/Q VGND VGND VPWR VPWR _19015_/Y sky130_fd_sc_hd__inv_2
X_16227_ _16227_/A VGND VGND VPWR VPWR _16227_/X sky130_fd_sc_hd__buf_2
XANTENNA__14184__A1 _14178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13439_ _13186_/Y _13431_/X _13438_/X VGND VGND VPWR VPWR _13439_/X sky130_fd_sc_hd__and3_4
XANTENNA__19647__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16158_ _16156_/Y _16154_/X _16157_/X _16154_/X VGND VGND VPWR VPWR _24694_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15109_ _24989_/Q _24593_/Q _15411_/A _15108_/Y VGND VGND VPWR VPWR _15116_/B sky130_fd_sc_hd__o22a_4
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16089_ _11730_/Y _15663_/X _15933_/X _24719_/Q _16088_/X VGND VGND VPWR VPWR _24719_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22799__A _22799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19917_ _19904_/Y VGND VGND VPWR VPWR _19917_/X sky130_fd_sc_hd__buf_2
XFILLER_142_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19848_ _23608_/Q VGND VGND VPWR VPWR _21763_/B sky130_fd_sc_hd__inv_2
XFILLER_69_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22311__B _22281_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16633__B1 _13599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19779_ _13403_/B VGND VGND VPWR VPWR _19779_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21810_ _21474_/A _20374_/Y VGND VGND VPWR VPWR _21812_/B sky130_fd_sc_hd__or2_4
XFILLER_25_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22790_ _22788_/X _22789_/X _22497_/X _16042_/A _22498_/X VGND VGND VPWR VPWR _22791_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17189__B2 _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21741_ _21741_/A _21740_/X VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__and2_4
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17421__A _14816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24460_ _25018_/CLK _16783_/X HRESETn VGND VGND VPWR VPWR _15022_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21672_ _21474_/A _21672_/B VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__or2_4
XFILLER_196_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _23555_/CLK _23411_/D VGND VGND VPWR VPWR _20383_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__20485__C _20499_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20623_ _20622_/Y VGND VGND VPWR VPWR _20623_/X sky130_fd_sc_hd__buf_2
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24391_ _24378_/CLK _24391_/D HRESETn VGND VGND VPWR VPWR _17045_/A sky130_fd_sc_hd__dfrtp_4
X_20554_ _20553_/X VGND VGND VPWR VPWR _23949_/D sky130_fd_sc_hd__inv_2
X_23342_ _16466_/A _23184_/X _21344_/X VGND VGND VPWR VPWR _23342_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24847__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15372__B1 _15348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20485_ _13893_/X _20682_/B _20499_/C VGND VGND VPWR VPWR _20486_/A sky130_fd_sc_hd__or3_4
X_23273_ _23273_/A VGND VGND VPWR VPWR _23273_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25012_ _25011_/CLK _25012_/D HRESETn VGND VGND VPWR VPWR _15321_/A sky130_fd_sc_hd__dfrtp_4
X_22224_ _22227_/A _19102_/Y VGND VGND VPWR VPWR _22224_/X sky130_fd_sc_hd__or2_4
XFILLER_180_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20799__A2 _20716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22155_ _24622_/Q _22155_/B VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__or2_4
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21106_ _24650_/Q _15663_/X _21105_/X _21049_/X VGND VGND VPWR VPWR _21106_/X sky130_fd_sc_hd__a211o_4
XFILLER_160_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_223_0_HCLK clkbuf_8_222_0_HCLK/A VGND VGND VPWR VPWR _25002_/CLK sky130_fd_sc_hd__clkbuf_1
X_22086_ _22394_/A _22086_/B VGND VGND VPWR VPWR _22087_/C sky130_fd_sc_hd__or2_4
XFILLER_248_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22502__A _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21037_ _21330_/A VGND VGND VPWR VPWR _22947_/A sky130_fd_sc_hd__buf_2
XFILLER_87_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16500__A _16495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16624__B1 _16364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12810_ _22724_/A VGND VGND VPWR VPWR _12858_/B sky130_fd_sc_hd__inv_2
XFILLER_228_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13790_ _13789_/X VGND VGND VPWR VPWR _21222_/B sky130_fd_sc_hd__inv_2
X_22988_ _23056_/A _22988_/B VGND VGND VPWR VPWR _22997_/C sky130_fd_sc_hd__and2_4
XANTENNA__22173__A1 _16532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12741_ _12739_/Y _12741_/B _12741_/C VGND VGND VPWR VPWR _25409_/D sky130_fd_sc_hd__and3_4
X_24727_ _24726_/CLK _24727_/D HRESETn VGND VGND VPWR VPWR _24727_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21939_ _21945_/A _21939_/B _21938_/X VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__and3_4
XFILLER_215_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17331__A _17331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15460_ _13963_/B _15458_/X _15455_/X _13963_/A _15453_/X VGND VGND VPWR VPWR _24971_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_179_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12672_ _12672_/A VGND VGND VPWR VPWR _25428_/D sky130_fd_sc_hd__inv_2
X_24658_ _24169_/CLK _24658_/D HRESETn VGND VGND VPWR VPWR _16263_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_179_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _20614_/A VGND VGND VPWR VPWR _20610_/A sky130_fd_sc_hd__inv_2
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23529_/CLK _23609_/D VGND VGND VPWR VPWR _23609_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _24994_/Q _15390_/Y VGND VGND VPWR VPWR _15391_/X sky130_fd_sc_hd__or2_4
XFILLER_179_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24589_ _24537_/CLK _16447_/X HRESETn VGND VGND VPWR VPWR _16445_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22891__B _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _17132_/B VGND VGND VPWR VPWR _17130_/Y sky130_fd_sc_hd__inv_2
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _12170_/X _14342_/B VGND VGND VPWR VPWR _14342_/X sky130_fd_sc_hd__or2_4
XFILLER_196_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24588__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17061_ _17062_/A _17062_/B VGND VGND VPWR VPWR _17061_/X sky130_fd_sc_hd__or2_4
X_14273_ _14268_/A VGND VGND VPWR VPWR _14273_/X sky130_fd_sc_hd__buf_2
XANTENNA__24517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16012_ _16019_/A VGND VGND VPWR VPWR _16012_/X sky130_fd_sc_hd__buf_2
X_13224_ _13217_/X _13220_/X _13223_/X VGND VGND VPWR VPWR _13224_/X sky130_fd_sc_hd__and3_4
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ _13212_/A VGND VGND VPWR VPWR _13155_/X sky130_fd_sc_hd__buf_2
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12106_ _12106_/A VGND VGND VPWR VPWR _12107_/A sky130_fd_sc_hd__buf_2
XANTENNA__16863__B1 _16726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13086_ _13006_/B _13080_/X _13083_/B _13040_/X VGND VGND VPWR VPWR _13087_/A sky130_fd_sc_hd__a211o_4
X_17963_ _17951_/A _17963_/B VGND VGND VPWR VPWR _17963_/X sky130_fd_sc_hd__or2_4
XFILLER_111_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22412__A _22854_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19702_ _19701_/Y _19699_/X _19656_/X _19699_/X VGND VGND VPWR VPWR _23659_/D sky130_fd_sc_hd__a2bb2o_4
X_12037_ _12036_/X VGND VGND VPWR VPWR _12050_/A sky130_fd_sc_hd__inv_2
X_16914_ _24281_/Q VGND VGND VPWR VPWR _16914_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17894_ _17896_/A _17891_/B _17894_/C VGND VGND VPWR VPWR _17894_/X sky130_fd_sc_hd__and3_4
XANTENNA__16410__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19633_ _19624_/Y VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__buf_2
XANTENNA__21028__A _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16845_ _16845_/A VGND VGND VPWR VPWR _16845_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16142__A1_N _16140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16776_ _16776_/A VGND VGND VPWR VPWR _16776_/Y sky130_fd_sc_hd__inv_2
X_19564_ _19564_/A VGND VGND VPWR VPWR _19564_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ _14011_/D VGND VGND VPWR VPWR _14027_/B sky130_fd_sc_hd__buf_2
XFILLER_230_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ _15726_/X VGND VGND VPWR VPWR _15727_/X sky130_fd_sc_hd__buf_2
X_18515_ _18515_/A _18515_/B _18486_/B _18473_/X VGND VGND VPWR VPWR _18516_/B sky130_fd_sc_hd__or4_4
XANTENNA__23243__A _23241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12939_ _12939_/A VGND VGND VPWR VPWR _25387_/D sky130_fd_sc_hd__inv_2
X_19495_ _23727_/Q VGND VGND VPWR VPWR _21691_/B sky130_fd_sc_hd__inv_2
XFILLER_207_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15658_ _16280_/A VGND VGND VPWR VPWR _15659_/B sky130_fd_sc_hd__buf_2
X_18446_ _16268_/Y _24167_/Q _23250_/A _18445_/Y VGND VGND VPWR VPWR _18451_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14609_ _14574_/X _14607_/Y _14608_/X _14599_/X _25094_/Q VGND VGND VPWR VPWR _14609_/X
+ sky130_fd_sc_hd__a32o_4
X_18377_ _18377_/A _25172_/Q _25167_/Q _14342_/B VGND VGND VPWR VPWR _18377_/X sky130_fd_sc_hd__or4_4
X_15589_ _15589_/A VGND VGND VPWR VPWR _15614_/A sky130_fd_sc_hd__buf_2
XFILLER_159_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17328_ _17263_/C _17332_/B _17327_/Y VGND VGND VPWR VPWR _17328_/X sky130_fd_sc_hd__o21a_4
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_231_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__24940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17259_ _17340_/A VGND VGND VPWR VPWR _17341_/A sky130_fd_sc_hd__inv_2
XFILLER_135_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19168__A _19181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20270_ _20270_/A VGND VGND VPWR VPWR _20270_/X sky130_fd_sc_hd__buf_2
XFILLER_190_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11729__A _14199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25248__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14105__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16854__B1 _16534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23960_ _23960_/CLK _20603_/X HRESETn VGND VGND VPWR VPWR _18887_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14759__B _14753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22911_ _22777_/X _22910_/X _22872_/X _24844_/Q _22779_/X VGND VGND VPWR VPWR _22911_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_53_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _24735_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_217_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23891_ _23889_/CLK _23891_/D VGND VGND VPWR VPWR _19034_/A sky130_fd_sc_hd__dfxtp_4
X_22842_ _15650_/X VGND VGND VPWR VPWR _22842_/X sky130_fd_sc_hd__buf_2
XANTENNA__21880__B _21867_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22773_ _12912_/A _22771_/X _22772_/X VGND VGND VPWR VPWR _22773_/X sky130_fd_sc_hd__o21a_4
X_24512_ _24509_/CLK _24512_/D HRESETn VGND VGND VPWR VPWR _16659_/A sky130_fd_sc_hd__dfrtp_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21724_ _21724_/A _21723_/X _21065_/X VGND VGND VPWR VPWR _21724_/X sky130_fd_sc_hd__or3_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25492_ _25494_/CLK _25492_/D HRESETn VGND VGND VPWR VPWR _12055_/A sky130_fd_sc_hd__dfrtp_4
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24443_ _24473_/CLK _16821_/X HRESETn VGND VGND VPWR VPWR _24443_/Q sky130_fd_sc_hd__dfrtp_4
X_21655_ _21217_/X VGND VGND VPWR VPWR _21972_/B sky130_fd_sc_hd__buf_2
XANTENNA__15593__B1 _11783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20606_ _20605_/X VGND VGND VPWR VPWR _20606_/Y sky130_fd_sc_hd__inv_2
X_24374_ _24639_/CLK _24374_/D HRESETn VGND VGND VPWR VPWR _24374_/Q sky130_fd_sc_hd__dfrtp_4
X_21586_ _21585_/X VGND VGND VPWR VPWR _21586_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24681__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23325_ _24648_/Q _21536_/X VGND VGND VPWR VPWR _23325_/X sky130_fd_sc_hd__or2_4
XFILLER_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20537_ _20537_/A _20537_/B VGND VGND VPWR VPWR _20543_/B sky130_fd_sc_hd__or2_4
XFILLER_153_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24610__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12159__B1 _12113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20468_ _24011_/Q _20456_/X _20461_/X _20469_/B VGND VGND VPWR VPWR _20468_/X sky130_fd_sc_hd__a211o_4
X_23256_ _14976_/A _22153_/X _22815_/X _23255_/X VGND VGND VPWR VPWR _23256_/X sky130_fd_sc_hd__a211o_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21969__A1 _21951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22207_ _22210_/A _22207_/B VGND VGND VPWR VPWR _22207_/X sky130_fd_sc_hd__or2_4
XFILLER_134_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19806__A _19788_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20399_ _21682_/B _20398_/X _19643_/A _20398_/X VGND VGND VPWR VPWR _20399_/X sky130_fd_sc_hd__a2bb2o_4
X_23187_ _23013_/A _23187_/B _23187_/C VGND VGND VPWR VPWR _23187_/X sky130_fd_sc_hd__and3_4
XANTENNA__20203__A2_N _20198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18710__A _18710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15648__B2 _15584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22138_ _21324_/X VGND VGND VPWR VPWR _22150_/A sky130_fd_sc_hd__buf_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14960_ _14960_/A _14960_/B _14957_/X _14959_/X VGND VGND VPWR VPWR _14993_/A sky130_fd_sc_hd__or4_4
XANTENNA__23040__C1 _23039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17326__A _17331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22069_ _22392_/A _19843_/Y VGND VGND VPWR VPWR _22071_/B sky130_fd_sc_hd__or2_4
X_13911_ _13963_/B VGND VGND VPWR VPWR _13911_/Y sky130_fd_sc_hd__inv_2
X_14891_ _14880_/X _14889_/Y _14837_/X _14890_/Y _14840_/A VGND VGND VPWR VPWR _14891_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16630_ _16629_/Y _16554_/A _16276_/X _16554_/A VGND VGND VPWR VPWR _16630_/X sky130_fd_sc_hd__a2bb2o_4
X_13842_ _13848_/A VGND VGND VPWR VPWR _13842_/X sky130_fd_sc_hd__buf_2
XFILLER_207_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23343__B1 _22852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16561_ _16558_/Y _16554_/X _16389_/X _16560_/X VGND VGND VPWR VPWR _24549_/D sky130_fd_sc_hd__a2bb2o_4
X_13773_ _13754_/X _13769_/X _13771_/X _14712_/A VGND VGND VPWR VPWR _25284_/D sky130_fd_sc_hd__o22a_4
X_15512_ _24947_/Q VGND VGND VPWR VPWR _15512_/Y sky130_fd_sc_hd__inv_2
X_18300_ _21212_/A _18300_/B VGND VGND VPWR VPWR _18301_/B sky130_fd_sc_hd__and2_4
X_12724_ _12728_/A _12718_/B _12724_/C VGND VGND VPWR VPWR _25415_/D sky130_fd_sc_hd__and3_4
X_19280_ _19280_/A VGND VGND VPWR VPWR _19280_/Y sky130_fd_sc_hd__inv_2
XFILLER_215_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16492_ _24574_/Q VGND VGND VPWR VPWR _16492_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24769__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18231_ _18231_/A _18231_/B VGND VGND VPWR VPWR _18233_/B sky130_fd_sc_hd__or2_4
X_15443_ _15443_/A VGND VGND VPWR VPWR _15447_/A sky130_fd_sc_hd__buf_2
X_12655_ _12636_/A _12655_/B _12655_/C VGND VGND VPWR VPWR _25433_/D sky130_fd_sc_hd__and3_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22449__A2 _22299_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ _18063_/A _18160_/X _18162_/C VGND VGND VPWR VPWR _18163_/C sky130_fd_sc_hd__and3_4
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _15380_/A _15384_/B VGND VGND VPWR VPWR _15381_/B sky130_fd_sc_hd__or2_4
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12618_/C _24875_/Q _12618_/C _24875_/Q VGND VGND VPWR VPWR _12586_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17113_ _16981_/Y _17117_/B _17112_/Y VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__o21a_4
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14315_/X _14324_/X _13493_/A _14320_/X VGND VGND VPWR VPWR _14325_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21311__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18093_ _18231_/A _18093_/B VGND VGND VPWR VPWR _18093_/X sky130_fd_sc_hd__or2_4
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17044_ _17105_/A _17016_/Y _17044_/C VGND VGND VPWR VPWR _17086_/D sky130_fd_sc_hd__or3_4
X_14256_ _13976_/A _14255_/X _13982_/A VGND VGND VPWR VPWR _14256_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19078__B2 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13207_ _13207_/A VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__buf_2
XANTENNA__17089__B1 _17065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14187_ _14174_/B _14181_/X _14182_/Y VGND VGND VPWR VPWR _14187_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_124_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22621__A2 _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13138_ _20725_/A _20725_/B _24024_/Q _20730_/A VGND VGND VPWR VPWR _13138_/X sky130_fd_sc_hd__or4_4
XANTENNA__25557__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18995_ _18994_/Y _18992_/X _18975_/X _18992_/X VGND VGND VPWR VPWR _23903_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22142__A _24489_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13069_ _13069_/A _13069_/B _13069_/C VGND VGND VPWR VPWR _13069_/X sky130_fd_sc_hd__and3_4
X_17946_ _17941_/X _17945_/X _18027_/A VGND VGND VPWR VPWR _17954_/B sky130_fd_sc_hd__o21a_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20396__B1 _19639_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17877_ _16901_/Y _17877_/B VGND VGND VPWR VPWR _17877_/X sky130_fd_sc_hd__or2_4
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19616_ _19614_/Y _19615_/X _19566_/X _19615_/X VGND VGND VPWR VPWR _23687_/D sky130_fd_sc_hd__a2bb2o_4
X_16828_ _16810_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__buf_2
XANTENNA__22137__A1 _13804_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19547_ _22404_/A VGND VGND VPWR VPWR _19547_/Y sky130_fd_sc_hd__inv_2
X_16759_ _15034_/Y _16758_/X _16410_/X _16758_/X VGND VGND VPWR VPWR _24472_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17013__B1 _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20699__B2 _20698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19478_ _19477_/Y _19473_/X _19410_/X _19460_/Y VGND VGND VPWR VPWR _23733_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18761__B1 _18714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18429_ _18429_/A _18424_/X _18429_/C _18429_/D VGND VGND VPWR VPWR _18430_/D sky130_fd_sc_hd__or4_4
XANTENNA__15575__B1 _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18108__A3 _18107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21440_ _21062_/A VGND VGND VPWR VPWR _21440_/X sky130_fd_sc_hd__buf_2
XFILLER_194_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21112__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21371_ _14885_/Y _21370_/X _14247_/Y _14230_/A VGND VGND VPWR VPWR _21377_/B sky130_fd_sc_hd__o22a_4
XFILLER_163_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16315__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20322_ _19527_/C _19986_/X _18289_/X VGND VGND VPWR VPWR _20323_/A sky130_fd_sc_hd__or3_4
X_23110_ _23110_/A VGND VGND VPWR VPWR _23110_/Y sky130_fd_sc_hd__inv_2
X_24090_ _24966_/CLK _24090_/D HRESETn VGND VGND VPWR VPWR _14290_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20253_ _20253_/A VGND VGND VPWR VPWR _20253_/Y sky130_fd_sc_hd__inv_2
X_23041_ _12268_/Y _22286_/X _22730_/X _12377_/Y _22858_/X VGND VGND VPWR VPWR _23041_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_162_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16827__B1 HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20184_ _20172_/A VGND VGND VPWR VPWR _20184_/X sky130_fd_sc_hd__buf_2
XANTENNA__23148__A _23148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24992_ _24966_/CLK _15406_/X HRESETn VGND VGND VPWR VPWR _15082_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23943_ _23395_/CLK _23943_/D HRESETn VGND VGND VPWR VPWR _23943_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23874_ _23871_/CLK _23874_/D VGND VGND VPWR VPWR _13270_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22128__A1 _21064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22825_ _22796_/X _22799_/X _22807_/Y _22824_/X VGND VGND VPWR VPWR HRDATA[16] sky130_fd_sc_hd__a211o_4
XANTENNA__16602__A1_N _16601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22679__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17004__B1 _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25544_ _24715_/CLK _11795_/X HRESETn VGND VGND VPWR VPWR _25544_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21887__B1 _24829_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22756_ _21058_/A _22755_/X _22303_/X _24875_/Q _22565_/X VGND VGND VPWR VPWR _22757_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_53_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24862__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21707_ _21700_/Y _21706_/Y _21526_/X VGND VGND VPWR VPWR _21707_/X sky130_fd_sc_hd__o21a_4
X_25475_ _23954_/CLK _25475_/D HRESETn VGND VGND VPWR VPWR _25475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_213_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22687_ _22687_/A VGND VGND VPWR VPWR _22687_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12440_ _12464_/A _12247_/X _12440_/C VGND VGND VPWR VPWR _12449_/D sky130_fd_sc_hd__or3_4
X_24426_ _24425_/CLK _24426_/D HRESETn VGND VGND VPWR VPWR _14931_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21638_ _21638_/A VGND VGND VPWR VPWR _22387_/A sky130_fd_sc_hd__buf_2
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13849__A _11851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _12370_/Y _24847_/Q _25350_/Q _12314_/Y VGND VGND VPWR VPWR _12380_/A sky130_fd_sc_hd__a2bb2o_4
X_24357_ _24625_/CLK _17363_/X HRESETn VGND VGND VPWR VPWR _24357_/Q sky130_fd_sc_hd__dfrtp_4
X_21569_ _21568_/Y _21161_/X _14877_/Y _21370_/X VGND VGND VPWR VPWR _21570_/A sky130_fd_sc_hd__o22a_4
XFILLER_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12753__A _25404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14110_ _14110_/A _14110_/B _14125_/A VGND VGND VPWR VPWR _14111_/B sky130_fd_sc_hd__or3_4
X_23308_ _23249_/A _23307_/X VGND VGND VPWR VPWR _23317_/B sky130_fd_sc_hd__nor2_4
XFILLER_154_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15090_ _15303_/A _24610_/Q _15303_/A _24610_/Q VGND VGND VPWR VPWR _15091_/D sky130_fd_sc_hd__a2bb2o_4
X_24288_ _25543_/CLK _24288_/D HRESETn VGND VGND VPWR VPWR _17752_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_176_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20142__A2_N _20141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14041_ _14032_/A VGND VGND VPWR VPWR _14043_/A sky130_fd_sc_hd__inv_2
XANTENNA__14541__A1 _25107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23239_ _23123_/X _23236_/Y _23168_/X _23238_/X VGND VGND VPWR VPWR _23239_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22603__A2 _23303_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17800_ _17798_/X _17800_/B _17799_/X VGND VGND VPWR VPWR _17801_/A sky130_fd_sc_hd__or3_4
X_15992_ _15797_/X _15895_/A _15775_/X _24757_/Q _15940_/X VGND VGND VPWR VPWR _15992_/X
+ sky130_fd_sc_hd__a32o_4
X_18780_ _18699_/B _18779_/X VGND VGND VPWR VPWR _18780_/X sky130_fd_sc_hd__or2_4
XFILLER_122_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22897__A _22897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14943_ _24428_/Q VGND VGND VPWR VPWR _14943_/Y sky130_fd_sc_hd__inv_2
X_17731_ _22266_/A VGND VGND VPWR VPWR _17732_/A sky130_fd_sc_hd__buf_2
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20378__B1 _19643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19271__A _19258_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14874_ _14832_/A _14822_/B _25049_/Q _14873_/X VGND VGND VPWR VPWR _14875_/A sky130_fd_sc_hd__a2bb2o_4
X_17662_ _17691_/A VGND VGND VPWR VPWR _17687_/A sky130_fd_sc_hd__buf_2
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19401_ _18111_/B VGND VGND VPWR VPWR _19401_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21590__A2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13825_ _13824_/X VGND VGND VPWR VPWR _21280_/A sky130_fd_sc_hd__inv_2
X_16613_ HWDATA[8] VGND VGND VPWR VPWR _16613_/X sky130_fd_sc_hd__buf_2
XANTENNA__21306__A _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17593_ _17610_/A _17610_/B VGND VGND VPWR VPWR _17594_/D sky130_fd_sc_hd__or2_4
XFILLER_223_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16544_ _24554_/Q VGND VGND VPWR VPWR _16544_/Y sky130_fd_sc_hd__inv_2
X_19332_ _19330_/Y _19325_/X _19308_/X _19331_/X VGND VGND VPWR VPWR _23786_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21878__B1 _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13756_ _13766_/A VGND VGND VPWR VPWR _13757_/C sky130_fd_sc_hd__buf_2
XFILLER_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12707_ _12728_/A _12705_/X _12706_/X VGND VGND VPWR VPWR _25419_/D sky130_fd_sc_hd__and3_4
X_16475_ _16540_/A VGND VGND VPWR VPWR _16495_/A sky130_fd_sc_hd__buf_2
X_19263_ _19263_/A VGND VGND VPWR VPWR _22070_/B sky130_fd_sc_hd__inv_2
X_13687_ _13686_/Y _11890_/X VGND VGND VPWR VPWR _13703_/B sky130_fd_sc_hd__or2_4
XANTENNA__24532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15426_ _15310_/A _15424_/X VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__or2_4
X_18214_ _17979_/A _18214_/B VGND VGND VPWR VPWR _18215_/C sky130_fd_sc_hd__or2_4
XFILLER_188_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12638_ _12702_/A _12638_/B VGND VGND VPWR VPWR _12647_/D sky130_fd_sc_hd__and2_4
X_19194_ _19193_/Y _19191_/X _19148_/X _19191_/X VGND VGND VPWR VPWR _23835_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15357_ _15357_/A _15357_/B _15356_/X VGND VGND VPWR VPWR _15358_/A sky130_fd_sc_hd__or3_4
X_18145_ _18039_/A _23783_/Q VGND VGND VPWR VPWR _18145_/X sky130_fd_sc_hd__or2_4
X_12569_ _25411_/Q VGND VGND VPWR VPWR _12713_/A sky130_fd_sc_hd__inv_2
XANTENNA__16135__A _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _14304_/A VGND VGND VPWR VPWR _14308_/Y sky130_fd_sc_hd__inv_2
X_18076_ _18039_/A _23785_/Q VGND VGND VPWR VPWR _18078_/B sky130_fd_sc_hd__or2_4
XFILLER_156_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15288_ _14990_/X _15291_/B _15183_/X VGND VGND VPWR VPWR _15288_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_116_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17027_ _17027_/A _17026_/X VGND VGND VPWR VPWR _17355_/B sky130_fd_sc_hd__or2_4
XFILLER_171_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14239_ _14237_/Y _14233_/X _13849_/X _14238_/X VGND VGND VPWR VPWR _14239_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15974__A _15796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16809__B1 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20605__A1 _14137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21802__B1 _13804_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18978_ _18977_/Y _18974_/X _18908_/X _18974_/X VGND VGND VPWR VPWR _18978_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17929_ _17929_/A VGND VGND VPWR VPWR _17929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19181__A _19181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20940_ _20944_/B _13674_/X VGND VGND VPWR VPWR _20940_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18982__B1 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20871_ _24055_/Q _20865_/X _20870_/X VGND VGND VPWR VPWR _20871_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_127_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _25030_/CLK sky130_fd_sc_hd__clkbuf_1
X_22610_ _24628_/Q _22610_/B VGND VGND VPWR VPWR _22610_/X sky130_fd_sc_hd__or2_4
XFILLER_223_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23590_ _23590_/CLK _23590_/D VGND VGND VPWR VPWR _19897_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22541_ _22541_/A VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__buf_2
XFILLER_195_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15548__B1 HADDR[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25260_ _25276_/CLK _25260_/D HRESETn VGND VGND VPWR VPWR _13857_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_50_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22472_ _22472_/A VGND VGND VPWR VPWR _22472_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14220__B1 _13812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24211_ _23522_/CLK _18348_/X HRESETn VGND VGND VPWR VPWR _13306_/A sky130_fd_sc_hd__dfrtp_4
X_21423_ _21387_/X _21388_/X _22523_/A _21422_/X VGND VGND VPWR VPWR _21423_/X sky130_fd_sc_hd__a211o_4
X_25191_ _25253_/CLK _25191_/D HRESETn VGND VGND VPWR VPWR _25191_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24142_ _24160_/CLK _24142_/D HRESETn VGND VGND VPWR VPWR _18604_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21354_ _21353_/X VGND VGND VPWR VPWR _21369_/B sky130_fd_sc_hd__inv_2
XANTENNA__25479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20305_ _20305_/A VGND VGND VPWR VPWR _22268_/B sky130_fd_sc_hd__inv_2
X_24073_ _24073_/CLK _24073_/D HRESETn VGND VGND VPWR VPWR _24073_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21285_ _25062_/Q _18277_/X VGND VGND VPWR VPWR _21285_/Y sky130_fd_sc_hd__nor2_4
XFILLER_104_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23024_ _16576_/A _22411_/X _15676_/X _23023_/X VGND VGND VPWR VPWR _23025_/C sky130_fd_sc_hd__a211o_4
X_20236_ _20232_/Y _20235_/X _19817_/X _20235_/X VGND VGND VPWR VPWR _23468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20167_ _20167_/A VGND VGND VPWR VPWR _21273_/B sky130_fd_sc_hd__inv_2
XANTENNA__25061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20098_ _20097_/Y _20093_/X _19761_/X _20093_/A VGND VGND VPWR VPWR _20098_/X sky130_fd_sc_hd__a2bb2o_4
X_24975_ _24975_/CLK _24975_/D HRESETn VGND VGND VPWR VPWR _13928_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22510__A _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19091__A _19091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11940_ _11938_/Y _11935_/X _11939_/X _11935_/X VGND VGND VPWR VPWR _11940_/X sky130_fd_sc_hd__a2bb2o_4
X_23926_ _23926_/CLK _23926_/D VGND VGND VPWR VPWR _18931_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_46_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_86_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_86_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11871_ _14248_/A VGND VGND VPWR VPWR _11871_/X sky130_fd_sc_hd__buf_2
X_23857_ _23871_/CLK _19129_/X VGND VGND VPWR VPWR _23857_/Q sky130_fd_sc_hd__dfxtp_4
X_13610_ _19054_/D VGND VGND VPWR VPWR _13610_/X sky130_fd_sc_hd__buf_2
X_22808_ _22808_/A VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__buf_2
XFILLER_32_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15124__A _15124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14590_ _14590_/A _14590_/B VGND VGND VPWR VPWR _14590_/X sky130_fd_sc_hd__or2_4
XFILLER_32_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23788_ _25082_/CLK _19327_/X VGND VGND VPWR VPWR _17958_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22521__A1 _13822_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13541_ _25309_/Q VGND VGND VPWR VPWR SSn_S2 sky130_fd_sc_hd__inv_2
X_25527_ _25528_/CLK _11868_/X HRESETn VGND VGND VPWR VPWR _25527_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23986__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22739_ _23010_/B VGND VGND VPWR VPWR _22827_/B sky130_fd_sc_hd__buf_2
XFILLER_241_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15539__B1 HADDR[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16260_ _16259_/Y _16257_/X _16157_/X _16257_/X VGND VGND VPWR VPWR _24660_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_197_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13472_ _13209_/A _13456_/X _13471_/X _25332_/Q _13208_/A VGND VGND VPWR VPWR _13472_/X
+ sky130_fd_sc_hd__o32a_4
X_25458_ _25456_/CLK _25458_/D HRESETn VGND VGND VPWR VPWR _25458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14211__B1 _13844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ _15201_/X VGND VGND VPWR VPWR _15215_/B sky130_fd_sc_hd__inv_2
X_12423_ _12261_/Y _12297_/X _12391_/X VGND VGND VPWR VPWR _12424_/B sky130_fd_sc_hd__or3_4
X_24409_ _24407_/CLK _24409_/D HRESETn VGND VGND VPWR VPWR _17062_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_200_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16191_ _16190_/X VGND VGND VPWR VPWR _16192_/A sky130_fd_sc_hd__buf_2
X_25389_ _25392_/CLK _25389_/D HRESETn VGND VGND VPWR VPWR _25389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15142_ _24994_/Q VGND VGND VPWR VPWR _15142_/Y sky130_fd_sc_hd__inv_2
X_12354_ _24830_/Q VGND VGND VPWR VPWR _12354_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15794__A _15793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22037__B1 _21697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15073_ _14930_/Y _15276_/A _15073_/C _15072_/X VGND VGND VPWR VPWR _15073_/X sky130_fd_sc_hd__or4_4
X_19950_ _23570_/Q VGND VGND VPWR VPWR _19950_/Y sky130_fd_sc_hd__inv_2
X_12285_ _25466_/Q VGND VGND VPWR VPWR _12401_/B sky130_fd_sc_hd__inv_2
XFILLER_5_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22404__B _21656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14024_ _13993_/X _14004_/X _14552_/A _14023_/X VGND VGND VPWR VPWR _14024_/X sky130_fd_sc_hd__a211o_4
X_18901_ _21002_/A VGND VGND VPWR VPWR _18901_/Y sky130_fd_sc_hd__inv_2
X_19881_ _19965_/A _18285_/D _19481_/X VGND VGND VPWR VPWR _19882_/A sky130_fd_sc_hd__or3_4
XFILLER_134_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12823__A1_N _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18832_ _16510_/Y _18657_/X _16510_/Y _18657_/X VGND VGND VPWR VPWR _18832_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11827__A _16252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14278__B1 _13809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18763_ _18763_/A _18751_/X VGND VGND VPWR VPWR _18764_/B sky130_fd_sc_hd__or2_4
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15975_ _15939_/X VGND VGND VPWR VPWR _15975_/X sky130_fd_sc_hd__buf_2
XANTENNA__22420__A _24624_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17714_ _17714_/A VGND VGND VPWR VPWR _21212_/A sky130_fd_sc_hd__buf_2
XFILLER_236_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14926_ _14924_/A _14925_/A _15016_/A _14925_/Y VGND VGND VPWR VPWR _14933_/B sky130_fd_sc_hd__o22a_4
X_18694_ _24146_/Q VGND VGND VPWR VPWR _18694_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24784__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18964__B1 _17430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _17577_/C _17644_/X VGND VGND VPWR VPWR _17646_/D sky130_fd_sc_hd__or2_4
XANTENNA__15778__B1 _24863_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14857_ _14854_/X _14856_/Y _25200_/Q _14854_/X VGND VGND VPWR VPWR _14857_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24713__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13808_ _25279_/Q VGND VGND VPWR VPWR _13808_/Y sky130_fd_sc_hd__inv_2
X_14788_ _14783_/A _14785_/X _14781_/X _14787_/Y VGND VGND VPWR VPWR _25064_/D sky130_fd_sc_hd__o22a_4
X_17576_ _24310_/Q VGND VGND VPWR VPWR _17644_/A sky130_fd_sc_hd__inv_2
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22512__A1 _14943_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19315_ _13396_/B VGND VGND VPWR VPWR _19315_/Y sky130_fd_sc_hd__inv_2
X_13739_ _13691_/X _13738_/Y _13689_/X _13722_/X _11702_/A VGND VGND VPWR VPWR _13739_/X
+ sky130_fd_sc_hd__a32o_4
X_16527_ _24560_/Q VGND VGND VPWR VPWR _16527_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19246_ _19131_/A VGND VGND VPWR VPWR _19246_/X sky130_fd_sc_hd__buf_2
X_16458_ _16192_/A VGND VGND VPWR VPWR _23009_/A sky130_fd_sc_hd__inv_2
X_15409_ _15120_/Y _15409_/B VGND VGND VPWR VPWR _15409_/Y sky130_fd_sc_hd__nand2_4
X_16389_ HWDATA[29] VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__buf_2
X_19177_ _19176_/Y _19174_/X _19085_/X _19174_/X VGND VGND VPWR VPWR _19177_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18128_ _18231_/A _18128_/B VGND VGND VPWR VPWR _18128_/X sky130_fd_sc_hd__or2_4
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18059_ _18059_/A VGND VGND VPWR VPWR _18138_/A sky130_fd_sc_hd__buf_2
XFILLER_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21070_ _15674_/A VGND VGND VPWR VPWR _21747_/A sky130_fd_sc_hd__buf_2
X_20021_ _20021_/A VGND VGND VPWR VPWR _20021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14269__B1 _13844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22968__C _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18645__A1_N _24537_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24760_ _24759_/CLK _15988_/X HRESETn VGND VGND VPWR VPWR _22418_/A sky130_fd_sc_hd__dfrtp_4
X_21972_ _19559_/Y _21972_/B VGND VGND VPWR VPWR _21972_/X sky130_fd_sc_hd__or2_4
XFILLER_67_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18955__B1 _18908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _23717_/CLK _23711_/D VGND VGND VPWR VPWR _23711_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _24067_/Q VGND VGND VPWR VPWR _20923_/Y sky130_fd_sc_hd__inv_2
XPHY_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24691_ _24689_/CLK _16165_/X HRESETn VGND VGND VPWR VPWR _22162_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15769__B1 _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _23642_/CLK _23642_/D VGND VGND VPWR VPWR _13297_/B sky130_fd_sc_hd__dfxtp_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ _20854_/A VGND VGND VPWR VPWR _20854_/X sky130_fd_sc_hd__buf_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _23493_/CLK _23573_/D VGND VGND VPWR VPWR _23573_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20785_ _20785_/A _20780_/Y VGND VGND VPWR VPWR _20785_/X sky130_fd_sc_hd__and2_4
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25312_ _25316_/CLK _25312_/D HRESETn VGND VGND VPWR VPWR _25312_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19380__B1 _19246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22524_ _13840_/Y _22524_/B VGND VGND VPWR VPWR _22524_/X sky130_fd_sc_hd__and2_4
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25243_ _25246_/CLK _14084_/X HRESETn VGND VGND VPWR VPWR _25243_/Q sky130_fd_sc_hd__dfrtp_4
X_22455_ _21449_/A VGND VGND VPWR VPWR _22487_/A sky130_fd_sc_hd__buf_2
XFILLER_167_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19132__B1 _19131_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21406_ _21262_/A _21396_/X _21405_/X VGND VGND VPWR VPWR _21406_/X sky130_fd_sc_hd__or3_4
XFILLER_136_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25174_ _24112_/CLK _14337_/X HRESETn VGND VGND VPWR VPWR _25174_/Q sky130_fd_sc_hd__dfrtp_4
X_22386_ _22090_/A _20057_/Y VGND VGND VPWR VPWR _22387_/C sky130_fd_sc_hd__or2_4
XFILLER_163_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24125_ _23946_/CLK _18898_/X HRESETn VGND VGND VPWR VPWR _24125_/Q sky130_fd_sc_hd__dfstp_4
X_21337_ _24420_/Q _21330_/X _21331_/X _21336_/X VGND VGND VPWR VPWR _21338_/C sky130_fd_sc_hd__a211o_4
XANTENNA__25242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12070_ _12070_/A VGND VGND VPWR VPWR _12070_/Y sky130_fd_sc_hd__inv_2
X_24056_ _24493_/CLK _24056_/D HRESETn VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21268_ _21638_/A _21266_/X _21267_/X VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__and3_4
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23007_ _20789_/Y _23006_/X _20928_/Y _21229_/X VGND VGND VPWR VPWR _23007_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17446__B1 _16729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20219_ _20213_/Y VGND VGND VPWR VPWR _20219_/X sky130_fd_sc_hd__buf_2
X_21199_ _24217_/Q _21199_/B VGND VGND VPWR VPWR _21199_/X sky130_fd_sc_hd__or2_4
XANTENNA__16938__A2_N _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15760_ _15758_/X _15751_/X _15759_/X _24872_/Q _15749_/X VGND VGND VPWR VPWR _15760_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_18_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17334__A _17212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12972_ _12969_/A _12969_/B VGND VGND VPWR VPWR _12972_/Y sky130_fd_sc_hd__nand2_4
X_24958_ _24138_/CLK _15487_/X HRESETn VGND VGND VPWR VPWR _24958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_92_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20348__A3 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18946__B1 _17433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ _11885_/X _11920_/Y VGND VGND VPWR VPWR _11923_/X sky130_fd_sc_hd__and2_4
X_14711_ _14709_/X _14710_/X _14709_/X _14710_/X VGND VGND VPWR VPWR _14711_/X sky130_fd_sc_hd__a2bb2o_4
X_15691_ _15696_/A _15696_/B _15691_/C VGND VGND VPWR VPWR _15691_/X sky130_fd_sc_hd__or3_4
X_23909_ _24111_/CLK _18980_/X VGND VGND VPWR VPWR _18979_/A sky130_fd_sc_hd__dfxtp_4
X_24889_ _24889_/CLK _15728_/X HRESETn VGND VGND VPWR VPWR _24889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12194__A1_N _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14642_ _14630_/X _14626_/Y _14641_/X _14624_/A _14631_/Y VGND VGND VPWR VPWR _25085_/D
+ sky130_fd_sc_hd__a32o_4
X_17430_ _14423_/A VGND VGND VPWR VPWR _17430_/X sky130_fd_sc_hd__buf_2
X_11854_ HWDATA[4] VGND VGND VPWR VPWR _11855_/A sky130_fd_sc_hd__buf_2
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20695__A _20716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_110_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24022_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _14610_/A _14610_/B VGND VGND VPWR VPWR _14574_/B sky130_fd_sc_hd__or2_4
X_17361_ _24357_/Q _17361_/B VGND VGND VPWR VPWR _17363_/B sky130_fd_sc_hd__or2_4
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ _25546_/Q VGND VGND VPWR VPWR _11785_/Y sky130_fd_sc_hd__inv_2
XFILLER_214_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_173_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23913_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19100_ _19099_/Y VGND VGND VPWR VPWR _19100_/X sky130_fd_sc_hd__buf_2
X_13524_ _14248_/A VGND VGND VPWR VPWR _13524_/X sky130_fd_sc_hd__buf_2
X_16312_ _16325_/A VGND VGND VPWR VPWR _16312_/X sky130_fd_sc_hd__buf_2
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17292_ _17294_/B VGND VGND VPWR VPWR _17292_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ _16240_/Y _16235_/X _16241_/X _16242_/X VGND VGND VPWR VPWR _16243_/X sky130_fd_sc_hd__a2bb2o_4
X_19031_ HWDATA[7] VGND VGND VPWR VPWR _19032_/A sky130_fd_sc_hd__buf_2
X_13455_ _13423_/A _13455_/B _13455_/C VGND VGND VPWR VPWR _13456_/C sky130_fd_sc_hd__or3_4
XFILLER_185_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ _12401_/B _12394_/D VGND VGND VPWR VPWR _12409_/B sky130_fd_sc_hd__or2_4
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16174_ _16173_/Y _16097_/X _15848_/X _16097_/X VGND VGND VPWR VPWR _24687_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ _13450_/A _18973_/A VGND VGND VPWR VPWR _13387_/C sky130_fd_sc_hd__or2_4
XANTENNA__17134__C1 _17065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12210__A2 _22871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15125_ _24983_/Q _15124_/A _15424_/A _15124_/Y VGND VGND VPWR VPWR _15125_/X sky130_fd_sc_hd__o22a_4
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12337_ _24854_/Q VGND VGND VPWR VPWR _12337_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12941__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15056_ _15056_/A _15052_/X _15054_/X _15055_/X VGND VGND VPWR VPWR _15056_/X sky130_fd_sc_hd__or4_4
X_19933_ _23577_/Q VGND VGND VPWR VPWR _19933_/Y sky130_fd_sc_hd__inv_2
X_12268_ _24775_/Q VGND VGND VPWR VPWR _12268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15160__B2 _24605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14007_ _13999_/B VGND VGND VPWR VPWR _14013_/B sky130_fd_sc_hd__buf_2
XANTENNA__17437__B1 _16791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19864_ _23603_/Q VGND VGND VPWR VPWR _22218_/B sky130_fd_sc_hd__inv_2
X_12199_ _22568_/A VGND VGND VPWR VPWR _12199_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18815_ _18809_/B VGND VGND VPWR VPWR _18815_/Y sky130_fd_sc_hd__inv_2
X_19795_ _19795_/A VGND VGND VPWR VPWR _22072_/B sky130_fd_sc_hd__inv_2
XFILLER_110_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18746_ _18733_/B _18710_/X _18733_/A VGND VGND VPWR VPWR _18746_/X sky130_fd_sc_hd__o21a_4
X_15958_ _12216_/Y _15953_/X _15957_/X _15953_/X VGND VGND VPWR VPWR _24777_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22733__B2 _22444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14909_ _14909_/A VGND VGND VPWR VPWR _14909_/Y sky130_fd_sc_hd__inv_2
X_18677_ _18749_/A VGND VGND VPWR VPWR _18739_/A sky130_fd_sc_hd__buf_2
X_15889_ _12831_/Y _15887_/X _11790_/X _15887_/X VGND VGND VPWR VPWR _24810_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17628_ _17621_/X VGND VGND VPWR VPWR _17629_/B sky130_fd_sc_hd__inv_2
XFILLER_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17559_ _11844_/Y _17504_/A _11859_/Y _24299_/Q VGND VGND VPWR VPWR _17560_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20570_ _20570_/A _20567_/A VGND VGND VPWR VPWR _20570_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16176__B1 _15489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19229_ _19228_/Y _19225_/X _19184_/X _19225_/X VGND VGND VPWR VPWR _19229_/X sky130_fd_sc_hd__a2bb2o_4
X_22240_ _22240_/A VGND VGND VPWR VPWR _22240_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22171_ _22171_/A _22171_/B _22171_/C VGND VGND VPWR VPWR _22171_/X sky130_fd_sc_hd__and3_4
XFILLER_173_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12851__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21122_ _21122_/A VGND VGND VPWR VPWR _21123_/A sky130_fd_sc_hd__buf_2
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17428__B1 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21053_ _21048_/X _21052_/Y _12989_/A _21048_/X VGND VGND VPWR VPWR _21053_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22421__B1 _16065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20004_ _21822_/B _19997_/X _20003_/X _19997_/X VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14778__A _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24635__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24812_ _24812_/CLK _15886_/X HRESETn VGND VGND VPWR VPWR _24812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24743_ _24372_/CLK _16029_/X HRESETn VGND VGND VPWR VPWR _16028_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_223_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21955_ _17727_/A _21955_/B VGND VGND VPWR VPWR _21957_/B sky130_fd_sc_hd__or2_4
XFILLER_55_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _24063_/Q VGND VGND VPWR VPWR _20906_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25135__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24674_ _24674_/CLK _16220_/X HRESETn VGND VGND VPWR VPWR _16219_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_70_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21886_ _16166_/Y _21436_/X _22662_/B _11853_/Y _21588_/X VGND VGND VPWR VPWR _21886_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15757__A3 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25198__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _23577_/CLK _23625_/D VGND VGND VPWR VPWR _23625_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _16728_/Y _20833_/X _24047_/Q _20836_/X VGND VGND VPWR VPWR _20837_/X sky130_fd_sc_hd__o22a_4
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23556_ _23555_/CLK _23556_/D VGND VGND VPWR VPWR _23556_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_246_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24966_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20768_ _20768_/A _20768_/B VGND VGND VPWR VPWR _20768_/X sky130_fd_sc_hd__or2_4
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22507_ _21542_/A VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__buf_2
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15914__B1 _24794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23494_/CLK _23487_/D VGND VGND VPWR VPWR _23487_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20699_ _15647_/Y _20695_/X _13131_/B _20698_/X VGND VGND VPWR VPWR _20699_/X sky130_fd_sc_hd__o22a_4
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _13285_/A _13225_/X _13240_/C VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__and3_4
X_25226_ _24095_/CLK _25226_/D HRESETn VGND VGND VPWR VPWR _25226_/Q sky130_fd_sc_hd__dfrtp_4
X_22438_ _22437_/X VGND VGND VPWR VPWR _22442_/A sky130_fd_sc_hd__buf_2
XFILLER_136_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14236__A1_N _14235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13171_ _13423_/A VGND VGND VPWR VPWR _13171_/X sky130_fd_sc_hd__buf_2
X_25157_ _24012_/CLK _14396_/X HRESETn VGND VGND VPWR VPWR _14395_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17329__A _17262_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22369_ _17732_/A _22368_/X _17738_/A VGND VGND VPWR VPWR _22369_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12761__A _25389_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12122_ _12122_/A VGND VGND VPWR VPWR _12122_/Y sky130_fd_sc_hd__inv_2
X_24108_ _23647_/CLK _24108_/D HRESETn VGND VGND VPWR VPWR _24108_/Q sky130_fd_sc_hd__dfrtp_4
X_25088_ _25276_/CLK _25088_/D HRESETn VGND VGND VPWR VPWR _13593_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12053_ _12052_/Y _12050_/X _25493_/Q _12050_/X VGND VGND VPWR VPWR _25494_/D sky130_fd_sc_hd__a2bb2o_4
X_16930_ _21531_/A _16929_/A _16171_/Y _16929_/Y VGND VGND VPWR VPWR _16931_/D sky130_fd_sc_hd__o22a_4
X_24039_ _24042_/CLK _24039_/D HRESETn VGND VGND VPWR VPWR _13145_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_151_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22963__B2 _22298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16861_ _19091_/A VGND VGND VPWR VPWR _16861_/X sky130_fd_sc_hd__buf_2
XANTENNA__24376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18600_ _24164_/Q _18599_/Y VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__or2_4
XANTENNA__16800__A2_N _16738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15812_ _12318_/Y _15808_/X _11766_/X _15811_/X VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17064__A _17064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19580_ _19574_/Y VGND VGND VPWR VPWR _19580_/X sky130_fd_sc_hd__buf_2
XFILLER_93_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16792_ _16737_/Y VGND VGND VPWR VPWR _16792_/X sky130_fd_sc_hd__buf_2
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18531_ _18531_/A _18531_/B VGND VGND VPWR VPWR _18534_/B sky130_fd_sc_hd__or2_4
XFILLER_46_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12955_ _12955_/A _12955_/B VGND VGND VPWR VPWR _12957_/B sky130_fd_sc_hd__or2_4
X_15743_ _12593_/Y _15741_/X _11790_/X _15741_/X VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_246_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17999__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18395__A1 _24121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11906_ _11905_/X _11898_/B VGND VGND VPWR VPWR _11906_/Y sky130_fd_sc_hd__nor2_4
X_18462_ _24193_/Q VGND VGND VPWR VPWR _18489_/A sky130_fd_sc_hd__inv_2
XFILLER_233_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12886_ _12638_/B _12863_/X VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__or2_4
X_15674_ _15674_/A VGND VGND VPWR VPWR _21574_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A VGND VGND VPWR VPWR _17413_/X sky130_fd_sc_hd__buf_2
XPHY_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _25533_/Q VGND VGND VPWR VPWR _11837_/Y sky130_fd_sc_hd__inv_2
X_14625_ _14624_/Y _13647_/A _14624_/A _13645_/X VGND VGND VPWR VPWR _14626_/B sky130_fd_sc_hd__o22a_4
X_18393_ _18393_/A VGND VGND VPWR VPWR _18393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12936__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19344__B1 _19254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11840__A _25532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14556_/A _14556_/B _14552_/X _14555_/X VGND VGND VPWR VPWR _14557_/A sky130_fd_sc_hd__or4_4
X_17344_ _17343_/X VGND VGND VPWR VPWR _24360_/D sky130_fd_sc_hd__inv_2
XANTENNA__16158__B1 _16157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11768_/A VGND VGND VPWR VPWR _11768_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21151__B1 _21577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _13516_/A VGND VGND VPWR VPWR _13507_/X sky130_fd_sc_hd__buf_2
XFILLER_202_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _14487_/A VGND VGND VPWR VPWR _14487_/Y sky130_fd_sc_hd__inv_2
X_17275_ _17242_/X _17272_/X _17274_/X VGND VGND VPWR VPWR _24377_/D sky130_fd_sc_hd__and3_4
XANTENNA__25164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11699_ _13690_/B _24231_/Q _13690_/B _24231_/Q VGND VGND VPWR VPWR _11699_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12719__B1 _12662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19014_ _19010_/Y _19004_/X _19012_/X _19013_/X VGND VGND VPWR VPWR _23898_/D sky130_fd_sc_hd__a2bb2o_4
X_13438_ _13332_/X _13434_/X _13438_/C VGND VGND VPWR VPWR _13438_/X sky130_fd_sc_hd__or3_4
X_16226_ _16226_/A VGND VGND VPWR VPWR _16226_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19127__A2_N _19121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22145__A _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16157_ HWDATA[8] VGND VGND VPWR VPWR _16157_/X sky130_fd_sc_hd__buf_2
X_13369_ _13369_/A _13369_/B VGND VGND VPWR VPWR _13370_/C sky130_fd_sc_hd__or2_4
XFILLER_155_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12671__A _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15108_ _24593_/Q VGND VGND VPWR VPWR _15108_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21984__A _19550_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16088_ _11729_/X _15668_/B VGND VGND VPWR VPWR _16088_/X sky130_fd_sc_hd__or2_4
XANTENNA__16330__B1 _15972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15133__B2 _15135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15039_ _24468_/Q VGND VGND VPWR VPWR _15039_/Y sky130_fd_sc_hd__inv_2
X_19916_ _23583_/Q VGND VGND VPWR VPWR _19916_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19454__A _19048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19847_ _21894_/B _19844_/X _19800_/X _19844_/X VGND VGND VPWR VPWR _23609_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19778_ _19777_/Y _19773_/X _19753_/X _19773_/X VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18729_ _18714_/A VGND VGND VPWR VPWR _18729_/X sky130_fd_sc_hd__buf_2
XFILLER_237_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16940__A1_N _16140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21740_ _16271_/Y _16192_/A _24588_/Q _16731_/Y VGND VGND VPWR VPWR _21740_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15739__A3 _15738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21671_ _21667_/X _21670_/X _17732_/X VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__o21a_4
XFILLER_196_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14947__B2 _14946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23410_ _23555_/CLK _23410_/D VGND VGND VPWR VPWR _20388_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11750__A _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20622_ _17411_/X VGND VGND VPWR VPWR _20622_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16955__A1_N _16169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ _24378_/CLK _17135_/Y HRESETn VGND VGND VPWR VPWR _24390_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16149__B1 _11827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21142__B1 _14191_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23341_ _23341_/A _22849_/X VGND VGND VPWR VPWR _23341_/X sky130_fd_sc_hd__or2_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20553_ _14178_/Y _20551_/X _20608_/A _20552_/X VGND VGND VPWR VPWR _20553_/X sky130_fd_sc_hd__a211o_4
XFILLER_177_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_13_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23565_/CLK sky130_fd_sc_hd__clkbuf_1
X_23272_ _21427_/A _23270_/X _22844_/X _23271_/X VGND VGND VPWR VPWR _23273_/A sky130_fd_sc_hd__o22a_4
XFILLER_164_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_76_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24759_/CLK sky130_fd_sc_hd__clkbuf_1
X_20484_ _25258_/Q _13871_/A _13862_/A VGND VGND VPWR VPWR _20499_/C sky130_fd_sc_hd__or3_4
XFILLER_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25011_ _25011_/CLK _25011_/D HRESETn VGND VGND VPWR VPWR _25011_/Q sky130_fd_sc_hd__dfrtp_4
X_22223_ _22210_/A _19283_/Y VGND VGND VPWR VPWR _22223_/X sky130_fd_sc_hd__or2_4
XFILLER_106_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22642__B1 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24887__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22154_ _21543_/A VGND VGND VPWR VPWR _22155_/B sky130_fd_sc_hd__buf_2
XANTENNA__22205__D _22204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16321__B1 _15963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24816__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21105_ _21021_/A _21105_/B VGND VGND VPWR VPWR _21105_/X sky130_fd_sc_hd__and2_4
XFILLER_121_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22085_ _22085_/A _22085_/B VGND VGND VPWR VPWR _22087_/B sky130_fd_sc_hd__or2_4
XFILLER_154_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22502__B _22662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21036_ _11744_/X VGND VGND VPWR VPWR _21330_/A sky130_fd_sc_hd__buf_2
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15978__A3 _16238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16908__A1_N _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22987_ _22488_/X _22985_/X _22986_/X _12535_/A _22784_/X VGND VGND VPWR VPWR _22988_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_216_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22173__A2 _21312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12740_ _12740_/A _12740_/B VGND VGND VPWR VPWR _12741_/B sky130_fd_sc_hd__or2_4
XFILLER_216_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21938_ _21938_/A _20046_/Y VGND VGND VPWR VPWR _21938_/X sky130_fd_sc_hd__or2_4
X_24726_ _24726_/CLK _16074_/X HRESETn VGND VGND VPWR VPWR _24726_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16388__B1 _16294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12671_ _12640_/B _12671_/B _12671_/C VGND VGND VPWR VPWR _12672_/A sky130_fd_sc_hd__or3_4
X_24657_ _24657_/CLK _16267_/X HRESETn VGND VGND VPWR VPWR _22107_/A sky130_fd_sc_hd__dfrtp_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _21330_/A VGND VGND VPWR VPWR _22424_/B sky130_fd_sc_hd__buf_2
XFILLER_188_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__A _12888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14408_/Y _14403_/X _14409_/X _14392_/X VGND VGND VPWR VPWR _25152_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _23513_/CLK _19849_/X VGND VGND VPWR VPWR _23608_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A VGND VGND VPWR VPWR _15390_/Y sky130_fd_sc_hd__inv_2
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _24523_/CLK _16449_/X HRESETn VGND VGND VPWR VPWR _24588_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _25173_/Q _14334_/X _14340_/Y VGND VGND VPWR VPWR _25173_/D sky130_fd_sc_hd__o21a_4
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ _23563_/CLK _23539_/D VGND VGND VPWR VPWR _23539_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _17060_/A _17059_/X VGND VGND VPWR VPWR _17062_/B sky130_fd_sc_hd__nor2_4
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _14272_/A VGND VGND VPWR VPWR _14272_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ _16004_/X VGND VGND VPWR VPWR _16019_/A sky130_fd_sc_hd__buf_2
X_13223_ _13222_/X _20260_/A VGND VGND VPWR VPWR _13223_/X sky130_fd_sc_hd__or2_4
X_25209_ _24523_/CLK _25209_/D HRESETn VGND VGND VPWR VPWR _14221_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17059__A _17074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13154_ _13153_/X VGND VGND VPWR VPWR _13177_/A sky130_fd_sc_hd__buf_2
XANTENNA__24557__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12105_ _17448_/A VGND VGND VPWR VPWR _12106_/A sky130_fd_sc_hd__buf_2
XFILLER_152_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13085_ _13104_/A _13085_/B _13085_/C VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__and3_4
X_17962_ _17943_/A _19412_/A VGND VGND VPWR VPWR _17962_/X sky130_fd_sc_hd__or2_4
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19701_ _23659_/Q VGND VGND VPWR VPWR _19701_/Y sky130_fd_sc_hd__inv_2
X_12036_ _25306_/Q _14299_/B _25311_/Q _25184_/Q VGND VGND VPWR VPWR _12036_/X sky130_fd_sc_hd__or4_4
X_16913_ _16913_/A _16913_/B _16911_/X _16912_/X VGND VGND VPWR VPWR _16932_/B sky130_fd_sc_hd__or4_4
X_17893_ _16936_/X _17858_/B VGND VGND VPWR VPWR _17894_/C sky130_fd_sc_hd__nand2_4
XFILLER_214_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19632_ _19632_/A VGND VGND VPWR VPWR _19632_/X sky130_fd_sc_hd__buf_2
XFILLER_238_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16844_ _16843_/Y _16839_/X _15759_/X _16839_/X VGND VGND VPWR VPWR _24431_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19563_ _19562_/Y _19557_/X _19402_/X _19557_/X VGND VGND VPWR VPWR _23704_/D sky130_fd_sc_hd__a2bb2o_4
X_16775_ _22682_/A _16773_/X _15756_/X _16773_/X VGND VGND VPWR VPWR _24464_/D sky130_fd_sc_hd__a2bb2o_4
X_13987_ _14027_/A VGND VGND VPWR VPWR _14053_/C sky130_fd_sc_hd__inv_2
X_18514_ _18514_/A VGND VGND VPWR VPWR _24189_/D sky130_fd_sc_hd__inv_2
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15726_ _15772_/A VGND VGND VPWR VPWR _15726_/X sky130_fd_sc_hd__buf_2
XFILLER_206_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12938_ _12912_/B _12911_/X _12883_/X _12934_/Y VGND VGND VPWR VPWR _12939_/A sky130_fd_sc_hd__a211o_4
X_19494_ _21825_/B _19489_/X _11957_/X _19489_/X VGND VGND VPWR VPWR _23728_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_230_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21044__A _24790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18445_ _24191_/Q VGND VGND VPWR VPWR _18445_/Y sky130_fd_sc_hd__inv_2
X_15657_ _15657_/A VGND VGND VPWR VPWR _16280_/A sky130_fd_sc_hd__buf_2
XANTENNA__25345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12869_ _12869_/A _12869_/B VGND VGND VPWR VPWR _12869_/X sky130_fd_sc_hd__or2_4
XPHY_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19317__B1 _19226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14608_ _14595_/A VGND VGND VPWR VPWR _14608_/X sky130_fd_sc_hd__buf_2
X_18376_ _18376_/A VGND VGND VPWR VPWR _18376_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15588_ _24921_/Q VGND VGND VPWR VPWR _15588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20883__A _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17327_ _17263_/C _17332_/B _17280_/X VGND VGND VPWR VPWR _17327_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14539_ _21352_/A _14519_/X _25107_/Q _14514_/X VGND VGND VPWR VPWR _14539_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17258_ _17258_/A VGND VGND VPWR VPWR _17258_/Y sky130_fd_sc_hd__inv_2
X_16209_ _23183_/A VGND VGND VPWR VPWR _16209_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17189_ _16374_/Y _17251_/A _16374_/Y _17251_/A VGND VGND VPWR VPWR _17190_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16303__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11729__B _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19184__A _19048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12876__C1 _12875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20938__B1 _20863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22910_ _22910_/A _23158_/B VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__or2_4
XANTENNA__15217__A _15293_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23890_ _23889_/CLK _19038_/X VGND VGND VPWR VPWR _23890_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22841_ _12255_/Y _23280_/A _22840_/X VGND VGND VPWR VPWR _22841_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_216_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23352__B2 _25062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22772_ _17766_/A _21457_/X _12464_/A _22447_/A VGND VGND VPWR VPWR _22772_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20166__B2 _20163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24511_ _24509_/CLK _24511_/D HRESETn VGND VGND VPWR VPWR _16662_/A sky130_fd_sc_hd__dfrtp_4
X_21723_ _17253_/Y _21321_/X _25376_/Q _21535_/A VGND VGND VPWR VPWR _21723_/X sky130_fd_sc_hd__a2bb2o_4
X_25491_ _25491_/CLK _12084_/X HRESETn VGND VGND VPWR VPWR _12072_/A sky130_fd_sc_hd__dfrtp_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16048__A _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24442_ _24473_/CLK _24442_/D HRESETn VGND VGND VPWR VPWR _16822_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21654_ _21384_/B VGND VGND VPWR VPWR _21654_/X sky130_fd_sc_hd__buf_2
XANTENNA__25015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20605_ _14137_/Y _20550_/Y _20564_/X _20604_/Y VGND VGND VPWR VPWR _20605_/X sky130_fd_sc_hd__a211o_4
X_24373_ _24372_/CLK _24373_/D HRESETn VGND VGND VPWR VPWR _17293_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22863__B1 _12568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21585_ _21578_/X _21581_/X _21582_/X _21584_/X VGND VGND VPWR VPWR _21585_/X sky130_fd_sc_hd__o22a_4
XFILLER_193_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23324_ _21714_/A _23324_/B VGND VGND VPWR VPWR _23331_/C sky130_fd_sc_hd__and2_4
X_20536_ _15465_/A _20521_/X _20534_/Y _20535_/X VGND VGND VPWR VPWR _20537_/B sky130_fd_sc_hd__a211o_4
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23255_ _24479_/Q _22673_/B _23190_/X VGND VGND VPWR VPWR _23255_/X sky130_fd_sc_hd__o21a_4
X_20467_ _14550_/A _20466_/Y VGND VGND VPWR VPWR _20469_/B sky130_fd_sc_hd__nor2_4
XFILLER_134_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21969__A2 _21966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22206_ _21398_/X VGND VGND VPWR VPWR _22210_/A sky130_fd_sc_hd__buf_2
X_23186_ _16566_/A _22940_/X _22941_/X _23185_/X VGND VGND VPWR VPWR _23187_/C sky130_fd_sc_hd__a211o_4
XFILLER_165_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20398_ _20385_/Y VGND VGND VPWR VPWR _20398_/X sky130_fd_sc_hd__buf_2
XFILLER_134_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22513__A _16524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24650__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22137_ _13804_/C _22101_/X _22105_/X _22111_/X _22136_/X VGND VGND VPWR VPWR _22137_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_161_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22918__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22068_ _21263_/A VGND VGND VPWR VPWR _22392_/A sky130_fd_sc_hd__buf_2
XFILLER_247_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12331__B2 _12330_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ _13910_/A VGND VGND VPWR VPWR _13963_/B sky130_fd_sc_hd__buf_2
X_21019_ sda_oen_o_S5 _24955_/Q _21012_/Y _15436_/A _21018_/Y VGND VGND VPWR VPWR
+ _23979_/D sky130_fd_sc_hd__a32o_4
XFILLER_102_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15127__A _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14890_ _24956_/Q VGND VGND VPWR VPWR _14890_/Y sky130_fd_sc_hd__inv_2
X_13841_ _13840_/Y _13838_/X _11834_/X _13838_/X VGND VGND VPWR VPWR _25269_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_242_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13772_ _13772_/A VGND VGND VPWR VPWR _14712_/A sky130_fd_sc_hd__buf_2
X_16560_ _16584_/A VGND VGND VPWR VPWR _16560_/X sky130_fd_sc_hd__buf_2
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20157__B2 _20156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15511_ _15510_/Y _15508_/X HADDR[18] _15508_/X VGND VGND VPWR VPWR _15511_/X sky130_fd_sc_hd__a2bb2o_4
X_12723_ _12621_/A _12723_/B VGND VGND VPWR VPWR _12724_/C sky130_fd_sc_hd__nand2_4
X_24709_ _24712_/CLK _24709_/D HRESETn VGND VGND VPWR VPWR _23061_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_204_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16491_ _16490_/Y _16488_/X _16315_/X _16488_/X VGND VGND VPWR VPWR _24575_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15033__B1 _25023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18230_ _18166_/A _18230_/B _18229_/X VGND VGND VPWR VPWR _18234_/B sky130_fd_sc_hd__and3_4
XFILLER_203_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15488__A1_N _14885_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12654_ _12642_/B _12654_/B VGND VGND VPWR VPWR _12655_/C sky130_fd_sc_hd__or2_4
X_15442_ _15439_/X VGND VGND VPWR VPWR _15443_/A sky130_fd_sc_hd__inv_2
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16781__B1 _11830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22449__A3 _22291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18161_ _18129_/A _19019_/A VGND VGND VPWR VPWR _18162_/C sky130_fd_sc_hd__or2_4
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15797__A _15796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _25421_/Q VGND VGND VPWR VPWR _12618_/C sky130_fd_sc_hd__inv_2
X_15373_ _15305_/A _15377_/B _15372_/Y VGND VGND VPWR VPWR _15373_/X sky130_fd_sc_hd__o21a_4
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21657__B2 _21656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _16981_/Y _17117_/B _17065_/X VGND VGND VPWR VPWR _17112_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ _25180_/Q _14311_/X _25179_/Q _14316_/X VGND VGND VPWR VPWR _14324_/X sky130_fd_sc_hd__o22a_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _18127_/A _18092_/B _18092_/C VGND VGND VPWR VPWR _18096_/B sky130_fd_sc_hd__and3_4
XFILLER_184_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24738__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14255_ _14255_/A _14255_/B VGND VGND VPWR VPWR _14255_/X sky130_fd_sc_hd__or2_4
X_17043_ _16996_/Y _17118_/A _17042_/X VGND VGND VPWR VPWR _17044_/C sky130_fd_sc_hd__or3_4
XANTENNA__22606__B1 _24871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ _13185_/X _13202_/X _13267_/A _25338_/Q _13207_/A VGND VGND VPWR VPWR _25338_/D
+ sky130_fd_sc_hd__a32o_4
X_14186_ _25136_/Q VGND VGND VPWR VPWR _14186_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13137_ _24021_/Q _13137_/B VGND VGND VPWR VPWR _20725_/B sky130_fd_sc_hd__or2_4
XANTENNA__12570__B2 _12572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18994_ _18994_/A VGND VGND VPWR VPWR _18994_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16421__A _24601_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22142__B _22854_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13068_ _13068_/A _13068_/B VGND VGND VPWR VPWR _13069_/C sky130_fd_sc_hd__nand2_4
X_17945_ _17945_/A _17945_/B _17945_/C VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__and3_4
XANTENNA__21039__A _22541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12019_ _12019_/A VGND VGND VPWR VPWR _12019_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17876_ _16937_/Y _17860_/D VGND VGND VPWR VPWR _17877_/B sky130_fd_sc_hd__or2_4
XFILLER_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20878__A _20836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19615_ _19615_/A VGND VGND VPWR VPWR _19615_/X sky130_fd_sc_hd__buf_2
X_16827_ _14978_/Y _16825_/X HWDATA[20] _16825_/X VGND VGND VPWR VPWR _24439_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22137__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23334__A1 _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17252__A _17362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19546_ _21192_/B _19541_/X _19501_/X _19528_/Y VGND VGND VPWR VPWR _23709_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12086__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16758_ _16762_/A VGND VGND VPWR VPWR _16758_/X sky130_fd_sc_hd__buf_2
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15709_ _16378_/A _16190_/B _16190_/C _15791_/D VGND VGND VPWR VPWR _15709_/X sky130_fd_sc_hd__or4_4
XFILLER_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17013__B2 _17050_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19477_ _19477_/A VGND VGND VPWR VPWR _19477_/Y sky130_fd_sc_hd__inv_2
X_16689_ _16689_/A VGND VGND VPWR VPWR _16689_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12396__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_26_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_26_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18428_ _16229_/A _24181_/Q _16229_/Y _18540_/A VGND VGND VPWR VPWR _18429_/D sky130_fd_sc_hd__o22a_4
XFILLER_221_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18359_ _18372_/A _18358_/X VGND VGND VPWR VPWR _18359_/Y sky130_fd_sc_hd__nand2_4
XFILLER_148_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18083__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15500__A _15503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21370_ _14443_/A VGND VGND VPWR VPWR _21370_/X sky130_fd_sc_hd__buf_2
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20321_ _23435_/Q VGND VGND VPWR VPWR _22365_/B sky130_fd_sc_hd__inv_2
XFILLER_163_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14116__A _14116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _22837_/X _23031_/Y _23035_/Y _23039_/X VGND VGND VPWR VPWR _23048_/C sky130_fd_sc_hd__a211o_4
X_20252_ _20251_/Y _20248_/X _19832_/X _20248_/X VGND VGND VPWR VPWR _20252_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20084__B1 _19769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17427__A _14420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20183_ _23487_/Q VGND VGND VPWR VPWR _20183_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14838__B1 _14235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16331__A _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24991_ _24975_/CLK _15408_/X HRESETn VGND VGND VPWR VPWR _24991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12313__B2 _24841_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19642__A _19624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23942_ _24095_/CLK _23942_/D HRESETn VGND VGND VPWR VPWR _22179_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23873_ _23871_/CLK _23873_/D VGND VGND VPWR VPWR _13307_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22128__A2 _22124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22824_ _22810_/Y _23020_/A _22824_/C _22824_/D VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__or4_4
XANTENNA__20139__B2 _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21887__A1 _24757_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22755_ _22755_/A _21104_/B VGND VGND VPWR VPWR _22755_/X sky130_fd_sc_hd__or2_4
X_25543_ _25543_/CLK _25543_/D HRESETn VGND VGND VPWR VPWR _25543_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21887__B2 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _21706_/A VGND VGND VPWR VPWR _21706_/Y sky130_fd_sc_hd__inv_2
X_25474_ _24119_/CLK _25474_/D HRESETn VGND VGND VPWR VPWR _12132_/A sky130_fd_sc_hd__dfrtp_4
X_22686_ _22459_/X _22683_/X _22462_/X _22685_/X VGND VGND VPWR VPWR _22687_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16763__B1 _16414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24425_ _24425_/CLK _16854_/X HRESETn VGND VGND VPWR VPWR _24425_/Q sky130_fd_sc_hd__dfrtp_4
X_21637_ _21611_/X _21637_/B _21636_/X VGND VGND VPWR VPWR _21637_/X sky130_fd_sc_hd__and3_4
XFILLER_200_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16506__A _16506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _12370_/A VGND VGND VPWR VPWR _12370_/Y sky130_fd_sc_hd__inv_2
X_24356_ _24354_/CLK _24356_/D HRESETn VGND VGND VPWR VPWR _17183_/A sky130_fd_sc_hd__dfrtp_4
X_21568_ _21568_/A VGND VGND VPWR VPWR _21568_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24831__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23307_ _20825_/Y _22298_/X _20964_/Y _22808_/X VGND VGND VPWR VPWR _23307_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20519_ _24089_/Q _20518_/X _14291_/X VGND VGND VPWR VPWR _20519_/X sky130_fd_sc_hd__o21a_4
X_24287_ _24272_/CLK _17810_/Y HRESETn VGND VGND VPWR VPWR _24287_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19817__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21499_ _22266_/A VGND VGND VPWR VPWR _21499_/X sky130_fd_sc_hd__buf_2
XFILLER_5_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23330__A1_N _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_46_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_46_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14040_ _14040_/A VGND VGND VPWR VPWR _14040_/Y sky130_fd_sc_hd__inv_2
X_23238_ _22563_/X _23237_/X _23062_/X _25553_/Q _23129_/X VGND VGND VPWR VPWR _23238_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_181_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22243__A _21210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13865__A _24007_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23169_ _22155_/B VGND VGND VPWR VPWR _23296_/B sky130_fd_sc_hd__buf_2
XANTENNA__16241__A _16241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23946__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15991_ _12241_/Y _15990_/X _15636_/X _15990_/X VGND VGND VPWR VPWR _15991_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13501__B1 _11871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12304__B2 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17730_ _17729_/Y VGND VGND VPWR VPWR _22266_/A sky130_fd_sc_hd__buf_2
X_14942_ _15072_/A VGND VGND VPWR VPWR _15271_/A sky130_fd_sc_hd__buf_2
XFILLER_209_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21575__B1 _15124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23074__A _23008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17661_ _17661_/A VGND VGND VPWR VPWR _17661_/Y sky130_fd_sc_hd__inv_2
X_14873_ _14873_/A _14873_/B _14889_/A _14832_/A VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__or4_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19400_ _19399_/Y _19397_/X _19377_/X _19397_/X VGND VGND VPWR VPWR _19400_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16612_ _16612_/A VGND VGND VPWR VPWR _16612_/Y sky130_fd_sc_hd__inv_2
X_13824_ _19595_/A _17422_/A VGND VGND VPWR VPWR _13824_/X sky130_fd_sc_hd__or2_4
X_17592_ _17571_/Y _17553_/Y _17573_/X _17591_/X VGND VGND VPWR VPWR _17610_/B sky130_fd_sc_hd__or4_4
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19331_ _19324_/Y VGND VGND VPWR VPWR _19331_/X sky130_fd_sc_hd__buf_2
X_16543_ _16542_/Y _16540_/X _16368_/X _16540_/X VGND VGND VPWR VPWR _16543_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11815__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21878__A1 _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13755_ _13754_/X VGND VGND VPWR VPWR _13772_/A sky130_fd_sc_hd__inv_2
XFILLER_231_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _12579_/Y _12704_/A VGND VGND VPWR VPWR _12706_/X sky130_fd_sc_hd__or2_4
X_19262_ _19261_/Y _19259_/X _16876_/X _19259_/X VGND VGND VPWR VPWR _23811_/D sky130_fd_sc_hd__a2bb2o_4
X_16474_ _16474_/A VGND VGND VPWR VPWR _16474_/Y sky130_fd_sc_hd__inv_2
X_13686_ _24225_/Q VGND VGND VPWR VPWR _13686_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _17977_/A _18213_/B VGND VGND VPWR VPWR _18213_/X sky130_fd_sc_hd__or2_4
X_15425_ _15310_/A _15424_/X VGND VGND VPWR VPWR _15425_/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12637_ _12730_/A VGND VGND VPWR VPWR _12640_/B sky130_fd_sc_hd__inv_2
X_19193_ _19193_/A VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__A _22678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18144_ _18037_/A _18142_/X _18143_/X VGND VGND VPWR VPWR _18144_/X sky130_fd_sc_hd__and3_4
X_12568_ _12568_/A VGND VGND VPWR VPWR _12568_/Y sky130_fd_sc_hd__inv_2
X_15356_ _15315_/X _15334_/D _15345_/C VGND VGND VPWR VPWR _15356_/X sky130_fd_sc_hd__o21a_4
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24572__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14307_ _14300_/A _14305_/X _14306_/Y VGND VGND VPWR VPWR _25186_/D sky130_fd_sc_hd__o21a_4
XFILLER_156_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18075_ _18037_/A _18073_/X _18074_/X VGND VGND VPWR VPWR _18075_/X sky130_fd_sc_hd__and3_4
X_12499_ _12218_/Y _12501_/B _12498_/Y VGND VGND VPWR VPWR _12499_/X sky130_fd_sc_hd__o21a_4
X_15287_ _15290_/A _15293_/B VGND VGND VPWR VPWR _15291_/B sky130_fd_sc_hd__or2_4
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17026_ _17007_/X _17026_/B _17026_/C _17025_/X VGND VGND VPWR VPWR _17026_/X sky130_fd_sc_hd__or4_4
XANTENNA__18259__B1 _17430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14238_ _14233_/A VGND VGND VPWR VPWR _14238_/X sky130_fd_sc_hd__buf_2
XANTENNA__23252__B1 _22852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22153__A _22947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16809__B2 _16806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14169_ _14169_/A VGND VGND VPWR VPWR _14169_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_3_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18977_ _23910_/Q VGND VGND VPWR VPWR _18977_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17928_ _13550_/A VGND VGND VPWR VPWR _17930_/A sky130_fd_sc_hd__inv_2
XFILLER_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17234__B2 _17391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17859_ _17757_/C _17858_/X VGND VGND VPWR VPWR _17860_/D sky130_fd_sc_hd__or2_4
XANTENNA__25360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15245__B1 _15208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23307__A1 _20825_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20870_ _20864_/Y _20859_/Y _20870_/C VGND VGND VPWR VPWR _20870_/X sky130_fd_sc_hd__and3_4
XFILLER_241_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21318__B1 _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19529_ _19528_/Y VGND VGND VPWR VPWR _19529_/X sky130_fd_sc_hd__buf_2
XFILLER_235_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11806__B1 _11805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22540_ _15095_/A _22589_/B VGND VGND VPWR VPWR _22548_/B sky130_fd_sc_hd__or2_4
XANTENNA__18860__A1_N _16517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15548__B2 _15547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22471_ _22468_/X _22469_/X _13822_/B _22470_/X VGND VGND VPWR VPWR _22472_/A sky130_fd_sc_hd__o22a_4
XFILLER_195_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22818__B1 _22815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24210_ _23522_/CLK _18350_/X HRESETn VGND VGND VPWR VPWR _13182_/A sky130_fd_sc_hd__dfrtp_4
X_21422_ _21180_/X _21406_/X _21421_/X VGND VGND VPWR VPWR _21422_/X sky130_fd_sc_hd__and3_4
X_25190_ _25253_/CLK _25190_/D HRESETn VGND VGND VPWR VPWR _14284_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24141_ _24160_/CLK _24141_/D HRESETn VGND VGND VPWR VPWR _24141_/Q sky130_fd_sc_hd__dfrtp_4
X_21353_ _21353_/A VGND VGND VPWR VPWR _21353_/X sky130_fd_sc_hd__buf_2
XFILLER_108_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20304_ _22344_/B _20303_/X _19990_/X _20303_/X VGND VGND VPWR VPWR _23443_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24072_ _24073_/CLK _20946_/X HRESETn VGND VGND VPWR VPWR _20944_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23159__A _22157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21284_ _21386_/B _21283_/X _13857_/Y _21386_/B VGND VGND VPWR VPWR _21284_/X sky130_fd_sc_hd__a2bb2o_4
X_23023_ _24574_/Q _22954_/B _22954_/C VGND VGND VPWR VPWR _23023_/X sky130_fd_sc_hd__and3_4
XFILLER_116_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20235_ _20234_/Y VGND VGND VPWR VPWR _20235_/X sky130_fd_sc_hd__buf_2
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20166_ _20165_/Y _20163_/X _20122_/X _20163_/X VGND VGND VPWR VPWR _20166_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15484__B1 _15483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20097_ _13453_/B VGND VGND VPWR VPWR _20097_/Y sky130_fd_sc_hd__inv_2
X_24974_ _24975_/CLK _15456_/X HRESETn VGND VGND VPWR VPWR _13929_/A sky130_fd_sc_hd__dfrtp_4
X_23925_ _23445_/CLK _23925_/D VGND VGND VPWR VPWR _18933_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11870_ HWDATA[1] VGND VGND VPWR VPWR _14248_/A sky130_fd_sc_hd__buf_2
XFILLER_217_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21126__B _21126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23856_ _23871_/CLK _19132_/X VGND VGND VPWR VPWR _19130_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_245_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16984__B1 _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22807_ _23072_/A _22807_/B VGND VGND VPWR VPWR _22807_/Y sky130_fd_sc_hd__nor2_4
X_20999_ _22179_/A _23943_/Q _21000_/B VGND VGND VPWR VPWR _23942_/D sky130_fd_sc_hd__o21a_4
X_23787_ _25082_/CLK _19329_/X VGND VGND VPWR VPWR _23787_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_213_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22521__A2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13540_ _20972_/B _13539_/X SCLK_S2 _20972_/B VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__a2bb2o_4
X_25526_ _24386_/CLK _25526_/D HRESETn VGND VGND VPWR VPWR _11869_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22738_ _22738_/A VGND VGND VPWR VPWR _23010_/B sky130_fd_sc_hd__buf_2
XANTENNA__15539__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13471_ _13186_/Y _13463_/X _13471_/C VGND VGND VPWR VPWR _13471_/X sky130_fd_sc_hd__and3_4
XFILLER_185_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22669_ _22669_/A _22669_/B VGND VGND VPWR VPWR _22669_/X sky130_fd_sc_hd__or2_4
X_25457_ _25456_/CLK _25457_/D HRESETn VGND VGND VPWR VPWR _25457_/Q sky130_fd_sc_hd__dfrtp_4
X_12422_ _12422_/A VGND VGND VPWR VPWR _25464_/D sky130_fd_sc_hd__inv_2
X_15210_ _15210_/A VGND VGND VPWR VPWR _15210_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24408_ _24407_/CLK _24408_/D HRESETn VGND VGND VPWR VPWR _24408_/Q sky130_fd_sc_hd__dfrtp_4
X_16190_ _16378_/A _16190_/B _16190_/C _16378_/D VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__or4_4
X_25388_ _25392_/CLK _25388_/D HRESETn VGND VGND VPWR VPWR _25388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _12353_/A VGND VGND VPWR VPWR _12353_/Y sky130_fd_sc_hd__inv_2
X_15141_ _15133_/X _15136_/X _15141_/C _15141_/D VGND VGND VPWR VPWR _15171_/A sky130_fd_sc_hd__or4_4
X_24339_ _24339_/CLK _17420_/X HRESETn VGND VGND VPWR VPWR _21018_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15072_ _15072_/A _15016_/A _15260_/C _15071_/X VGND VGND VPWR VPWR _15072_/X sky130_fd_sc_hd__or4_4
XFILLER_5_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20357__A1_N _20356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12284_ _12514_/A VGND VGND VPWR VPWR _12398_/A sky130_fd_sc_hd__buf_2
XANTENNA__23069__A _16671_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14023_ _14553_/A _14556_/A _14553_/A _14556_/A VGND VGND VPWR VPWR _14023_/X sky130_fd_sc_hd__a2bb2o_4
X_18900_ _24013_/Q _14544_/Y _21000_/A _14543_/A VGND VGND VPWR VPWR _18900_/X sky130_fd_sc_hd__o22a_4
X_19880_ _23596_/Q VGND VGND VPWR VPWR _22346_/B sky130_fd_sc_hd__inv_2
X_18831_ _16502_/Y _24149_/Q _16502_/Y _24149_/Q VGND VGND VPWR VPWR _18831_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_133_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _24206_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_1_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15475__B1 _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_196_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24488_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15102__A2_N _24585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18762_ _18698_/C _18766_/B _18761_/Y VGND VGND VPWR VPWR _18762_/X sky130_fd_sc_hd__o21a_4
X_15974_ _15796_/X VGND VGND VPWR VPWR _15974_/X sky130_fd_sc_hd__buf_2
XANTENNA__25118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22420__B _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17713_ _17898_/B VGND VGND VPWR VPWR _17713_/X sky130_fd_sc_hd__buf_2
XFILLER_208_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14925_ _14925_/A VGND VGND VPWR VPWR _14925_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21317__A _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18693_ _18693_/A VGND VGND VPWR VPWR _18699_/B sky130_fd_sc_hd__inv_2
XFILLER_209_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17644_ _17644_/A _17635_/X VGND VGND VPWR VPWR _17644_/X sky130_fd_sc_hd__or2_4
X_14856_ _14856_/A VGND VGND VPWR VPWR _14856_/Y sky130_fd_sc_hd__inv_2
X_13807_ _13795_/Y _13805_/X _13806_/X _13805_/X VGND VGND VPWR VPWR _13807_/X sky130_fd_sc_hd__a2bb2o_4
X_17575_ _17575_/A VGND VGND VPWR VPWR _17577_/C sky130_fd_sc_hd__inv_2
XFILLER_189_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14787_ _14787_/A VGND VGND VPWR VPWR _14787_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16663__A1_N _16662_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11999_ _25319_/Q VGND VGND VPWR VPWR _11999_/Y sky130_fd_sc_hd__inv_2
X_19314_ _19313_/Y _19309_/X _19246_/X _19309_/X VGND VGND VPWR VPWR _19314_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16526_ _16524_/Y _16520_/X _16153_/X _16525_/X VGND VGND VPWR VPWR _16526_/X sky130_fd_sc_hd__a2bb2o_4
X_13738_ _13691_/A _13690_/X VGND VGND VPWR VPWR _13738_/Y sky130_fd_sc_hd__nand2_4
XFILLER_177_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16727__B1 _16726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22148__A _21607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24753__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19245_ _13349_/B VGND VGND VPWR VPWR _19245_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16457_ _18515_/A VGND VGND VPWR VPWR _18488_/A sky130_fd_sc_hd__buf_2
X_13669_ _24057_/Q _13668_/X VGND VGND VPWR VPWR _13670_/B sky130_fd_sc_hd__or2_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15408_ _15393_/A _15408_/B _15408_/C VGND VGND VPWR VPWR _15408_/X sky130_fd_sc_hd__and3_4
X_19176_ _18100_/B VGND VGND VPWR VPWR _19176_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25310__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16388_ _16387_/Y _16384_/X _16294_/X _16384_/X VGND VGND VPWR VPWR _24615_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12393__B _13017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18127_ _18127_/A _18125_/X _18127_/C VGND VGND VPWR VPWR _18131_/B sky130_fd_sc_hd__and3_4
X_15339_ _25008_/Q _15343_/B VGND VGND VPWR VPWR _15341_/B sky130_fd_sc_hd__or2_4
XFILLER_172_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18058_ _18131_/A _18054_/X _18057_/X VGND VGND VPWR VPWR _18069_/B sky130_fd_sc_hd__or3_4
XFILLER_144_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17009_ _16026_/Y _24401_/Q _16026_/Y _24401_/Q VGND VGND VPWR VPWR _17012_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_92_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_92_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20020_ _20019_/Y _20017_/X _19993_/X _20017_/X VGND VGND VPWR VPWR _23547_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21539__B1 _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17207__A1 _24626_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17207__B2 _17364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21971_ _21971_/A _21971_/B VGND VGND VPWR VPWR _21971_/X sky130_fd_sc_hd__or2_4
XFILLER_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12849__A _25401_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20922_ _20921_/X VGND VGND VPWR VPWR _24066_/D sky130_fd_sc_hd__inv_2
X_23710_ _23717_/CLK _23710_/D VGND VGND VPWR VPWR _23710_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24690_ _24689_/CLK _16168_/X HRESETn VGND VGND VPWR VPWR _16166_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20853_ _20852_/X VGND VGND VPWR VPWR _20853_/Y sky130_fd_sc_hd__inv_2
X_23641_ _23631_/CLK _19751_/X VGND VGND VPWR VPWR _19750_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_199_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23513_/CLK _23572_/D VGND VGND VPWR VPWR _19944_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20784_ _20790_/B VGND VGND VPWR VPWR _20785_/A sky130_fd_sc_hd__inv_2
XANTENNA__24494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _22523_/A VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__buf_2
X_25311_ _25188_/CLK _25311_/D HRESETn VGND VGND VPWR VPWR _25311_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22454_ _17861_/B _22446_/A _25381_/Q _22453_/X VGND VGND VPWR VPWR _22454_/X sky130_fd_sc_hd__a2bb2o_4
X_25242_ _25246_/CLK _25242_/D HRESETn VGND VGND VPWR VPWR _13999_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_194_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21405_ _21401_/X _21404_/X _25068_/Q VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__o21a_4
X_25173_ _24112_/CLK _25173_/D HRESETn VGND VGND VPWR VPWR _25173_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15895__A _15895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22385_ _22385_/A _22385_/B VGND VGND VPWR VPWR _22387_/B sky130_fd_sc_hd__or2_4
XFILLER_194_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24124_ _23946_/CLK _18899_/X HRESETn VGND VGND VPWR VPWR _24124_/Q sky130_fd_sc_hd__dfstp_4
X_21336_ _24452_/Q _21312_/B _21335_/X VGND VGND VPWR VPWR _21336_/X sky130_fd_sc_hd__o21a_4
XFILLER_136_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24055_ _24493_/CLK _24055_/D HRESETn VGND VGND VPWR VPWR _24055_/Q sky130_fd_sc_hd__dfrtp_4
X_21267_ _21267_/A _20209_/Y VGND VGND VPWR VPWR _21267_/X sky130_fd_sc_hd__or2_4
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23006_ _21123_/X VGND VGND VPWR VPWR _23006_/X sky130_fd_sc_hd__buf_2
X_20218_ _23474_/Q VGND VGND VPWR VPWR _20218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21198_ _18319_/A _21189_/X _21197_/X VGND VGND VPWR VPWR _21198_/X sky130_fd_sc_hd__or3_4
Xclkbuf_8_206_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _24523_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20149_ _19859_/X _20149_/B _18914_/X VGND VGND VPWR VPWR _20149_/X sky130_fd_sc_hd__or3_4
XFILLER_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23336__B _16552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21137__A _25107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12971_ _12783_/Y _12969_/X _12970_/Y VGND VGND VPWR VPWR _25380_/D sky130_fd_sc_hd__o21a_4
X_24957_ _24138_/CLK _24957_/D HRESETn VGND VGND VPWR VPWR _14885_/A sky130_fd_sc_hd__dfstp_4
XFILLER_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15209__B1 _15208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14710_ _13762_/X _14693_/A _13744_/X _14693_/Y VGND VGND VPWR VPWR _14710_/X sky130_fd_sc_hd__o22a_4
XFILLER_245_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21545__A3 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15135__A _15135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11922_ _11879_/A _11893_/X _11920_/Y _11887_/A _11921_/Y VGND VGND VPWR VPWR _25519_/D
+ sky130_fd_sc_hd__a32o_4
X_23908_ _23885_/CLK _23908_/D VGND VGND VPWR VPWR _18981_/A sky130_fd_sc_hd__dfxtp_4
X_15690_ _24892_/Q VGND VGND VPWR VPWR _15696_/B sky130_fd_sc_hd__inv_2
XFILLER_206_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24888_ _24889_/CLK _24888_/D HRESETn VGND VGND VPWR VPWR _12591_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14641_ _14626_/A _14626_/B VGND VGND VPWR VPWR _14641_/X sky130_fd_sc_hd__or2_4
X_11853_ _11853_/A VGND VGND VPWR VPWR _11853_/Y sky130_fd_sc_hd__inv_2
X_23839_ _24101_/CLK _19182_/X VGND VGND VPWR VPWR _19180_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _17360_/A VGND VGND VPWR VPWR _17361_/B sky130_fd_sc_hd__inv_2
XFILLER_198_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _11782_/Y _11777_/X _11783_/X _11777_/X VGND VGND VPWR VPWR _25547_/D sky130_fd_sc_hd__a2bb2o_4
X_14572_ _14613_/A _14613_/B VGND VGND VPWR VPWR _14610_/B sky130_fd_sc_hd__or2_4
XFILLER_202_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _23091_/A VGND VGND VPWR VPWR _16311_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ _13523_/A VGND VGND VPWR VPWR _13536_/A sky130_fd_sc_hd__inv_2
X_25509_ _23678_/CLK _25509_/D HRESETn VGND VGND VPWR VPWR _20010_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17291_ _17345_/A _17267_/X VGND VGND VPWR VPWR _17294_/B sky130_fd_sc_hd__or2_4
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19030_ _19037_/A VGND VGND VPWR VPWR _19030_/X sky130_fd_sc_hd__buf_2
X_16242_ _16264_/A VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__buf_2
X_13454_ _13454_/A _13454_/B _13454_/C VGND VGND VPWR VPWR _13455_/C sky130_fd_sc_hd__and3_4
X_12405_ _12405_/A VGND VGND VPWR VPWR _12405_/Y sky130_fd_sc_hd__inv_2
X_13385_ _13385_/A _13385_/B VGND VGND VPWR VPWR _13385_/X sky130_fd_sc_hd__or2_4
X_16173_ _21444_/A VGND VGND VPWR VPWR _16173_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15124_ _15124_/A VGND VGND VPWR VPWR _15124_/Y sky130_fd_sc_hd__inv_2
X_12336_ _13023_/A VGND VGND VPWR VPWR _13024_/A sky130_fd_sc_hd__inv_2
XFILLER_154_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11838__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_16_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_12267_ _12299_/A _24779_/Q _25458_/Q _12266_/Y VGND VGND VPWR VPWR _12267_/X sky130_fd_sc_hd__a2bb2o_4
X_15055_ _14912_/X _15034_/Y _15195_/A _15024_/Y VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__a2bb2o_4
X_19932_ _22094_/B _19926_/X _19796_/X _19931_/X VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21769__B1 _14721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14006_ _13999_/A VGND VGND VPWR VPWR _14013_/A sky130_fd_sc_hd__buf_2
X_19863_ _19858_/Y _19862_/X _19790_/X _19862_/X VGND VGND VPWR VPWR _19863_/X sky130_fd_sc_hd__a2bb2o_4
X_12198_ _12197_/X _22778_/A _12197_/A _22778_/A VGND VGND VPWR VPWR _12198_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22431__A _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18814_ _18806_/A _18810_/X _18813_/Y VGND VGND VPWR VPWR _24137_/D sky130_fd_sc_hd__and3_4
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19794_ _22233_/B _19789_/X _19793_/X _19789_/X VGND VGND VPWR VPWR _23627_/D sky130_fd_sc_hd__a2bb2o_4
X_18745_ _18739_/A _18735_/B _18745_/C VGND VGND VPWR VPWR _18745_/X sky130_fd_sc_hd__and3_4
XANTENNA__21047__A _21046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15957_ HWDATA[24] VGND VGND VPWR VPWR _15957_/X sky130_fd_sc_hd__buf_2
XFILLER_110_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14908_ _15231_/A _24435_/Q _14906_/Y _24435_/Q VGND VGND VPWR VPWR _14919_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18676_ _18713_/A VGND VGND VPWR VPWR _18749_/A sky130_fd_sc_hd__buf_2
X_15888_ _12767_/Y _15887_/X _11787_/X _15887_/X VGND VGND VPWR VPWR _15888_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17627_ _17598_/A _17627_/B _17626_/Y VGND VGND VPWR VPWR _17627_/X sky130_fd_sc_hd__and3_4
XFILLER_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14839_ _14834_/X _14838_/X _14806_/A _14834_/X VGND VGND VPWR VPWR _25060_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17558_ _25553_/Q _17569_/A _11853_/Y _24300_/Q VGND VGND VPWR VPWR _17558_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16509_ _16506_/Y _16508_/X _16334_/X _16508_/X VGND VGND VPWR VPWR _16509_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17489_ _11661_/A _17484_/X _18361_/A VGND VGND VPWR VPWR _24329_/D sky130_fd_sc_hd__a21oi_4
X_19228_ _23822_/Q VGND VGND VPWR VPWR _19228_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19159_ _19159_/A VGND VGND VPWR VPWR _19159_/X sky130_fd_sc_hd__buf_2
XANTENNA__16604__A _16618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22170_ _24425_/Q _21330_/X _21331_/X _22169_/X VGND VGND VPWR VPWR _22171_/C sky130_fd_sc_hd__a211o_4
XFILLER_133_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12851__B _12952_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21121_ _21121_/A VGND VGND VPWR VPWR _21121_/X sky130_fd_sc_hd__buf_2
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21052_ _21051_/X VGND VGND VPWR VPWR _21052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22421__A1 _22289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22421__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16555__A1_N _16550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20003_ _20003_/A VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__buf_2
XFILLER_219_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24811_ _24856_/CLK _15888_/X HRESETn VGND VGND VPWR VPWR _22985_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20499__C _20499_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_36_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _23926_/CLK sky130_fd_sc_hd__clkbuf_1
X_24742_ _24642_/CLK _24742_/D HRESETn VGND VGND VPWR VPWR _24742_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21954_ _17716_/A _21952_/X _21953_/X VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__and3_4
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_99_0_HCLK clkbuf_7_49_0_HCLK/X VGND VGND VPWR VPWR _24651_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24675__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20905_ _20900_/X _20903_/Y _24499_/Q _20904_/X VGND VGND VPWR VPWR _20905_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_243_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21103_/A VGND VGND VPWR VPWR _22662_/B sky130_fd_sc_hd__buf_2
X_24673_ _24552_/CLK _16223_/X HRESETn VGND VGND VPWR VPWR _24673_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24604__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20836_/A VGND VGND VPWR VPWR _20836_/X sky130_fd_sc_hd__buf_2
X_23624_ _23529_/CLK _23624_/D VGND VGND VPWR VPWR _19802_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_187_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _20768_/A VGND VGND VPWR VPWR _20772_/A sky130_fd_sc_hd__inv_2
X_23555_ _23555_/CLK _23555_/D VGND VGND VPWR VPWR _23555_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _22436_/X _22487_/X _22506_/C _22505_/X VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__or4_4
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23486_ _23494_/CLK _20187_/X VGND VGND VPWR VPWR _23486_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20698_ _20788_/A VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__buf_2
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22516__A _21596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22437_ _21321_/A VGND VGND VPWR VPWR _22437_/X sky130_fd_sc_hd__buf_2
X_25225_ _23395_/CLK _14154_/X HRESETn VGND VGND VPWR VPWR _14111_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_136_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13170_ _13182_/A VGND VGND VPWR VPWR _13423_/A sky130_fd_sc_hd__inv_2
X_22368_ _17716_/A _22364_/X _22365_/X _22366_/X _22367_/X VGND VGND VPWR VPWR _22368_/X
+ sky130_fd_sc_hd__a32o_4
X_25156_ _24012_/CLK _14398_/X HRESETn VGND VGND VPWR VPWR _20438_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18864__B1 _16512_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12121_ _12120_/Y _12116_/X _11851_/X _12116_/X VGND VGND VPWR VPWR _25479_/D sky130_fd_sc_hd__a2bb2o_4
X_21319_ _22723_/A _21318_/X VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__and2_4
X_24107_ _23647_/CLK _24107_/D HRESETn VGND VGND VPWR VPWR _24107_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22323__A1_N _14116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25087_ _23703_/CLK _25087_/D HRESETn VGND VGND VPWR VPWR _25087_/Q sky130_fd_sc_hd__dfrtp_4
X_22299_ _15631_/Y _22299_/B VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__and2_4
XFILLER_124_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ _25494_/Q VGND VGND VPWR VPWR _12052_/Y sky130_fd_sc_hd__inv_2
X_24038_ _24500_/CLK _24038_/D HRESETn VGND VGND VPWR VPWR _20797_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17419__B2 _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16860_ _16859_/Y _16857_/X _16796_/X _16857_/X VGND VGND VPWR VPWR _24422_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17345__A _17345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15811_ _15818_/A VGND VGND VPWR VPWR _15811_/X sky130_fd_sc_hd__buf_2
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22401__D _22401_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16791_ _19085_/A VGND VGND VPWR VPWR _16791_/X sky130_fd_sc_hd__buf_2
XFILLER_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18530_ _18472_/X _18538_/B VGND VGND VPWR VPWR _18531_/B sky130_fd_sc_hd__or2_4
XFILLER_219_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15850__B1 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ _12535_/Y _15741_/X _11787_/X _15741_/X VGND VGND VPWR VPWR _24881_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19560__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ _12956_/B VGND VGND VPWR VPWR _12955_/B sky130_fd_sc_hd__inv_2
XFILLER_246_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18395__A2 _18377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11905_ _17711_/A VGND VGND VPWR VPWR _11905_/X sky130_fd_sc_hd__buf_2
X_18461_ _18493_/A VGND VGND VPWR VPWR _18492_/A sky130_fd_sc_hd__buf_2
X_15673_ _15673_/A VGND VGND VPWR VPWR _15674_/A sky130_fd_sc_hd__buf_2
XFILLER_206_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12885_ _12885_/A VGND VGND VPWR VPWR _25401_/D sky130_fd_sc_hd__inv_2
Xclkbuf_5_7_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17411_/X VGND VGND VPWR VPWR _17413_/A sky130_fd_sc_hd__buf_2
X_14624_ _14624_/A VGND VGND VPWR VPWR _14624_/Y sky130_fd_sc_hd__inv_2
XPHY_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11833_/Y _11825_/X _11834_/X _11835_/X VGND VGND VPWR VPWR _25534_/D sky130_fd_sc_hd__a2bb2o_4
X_18392_ _18390_/Y _18391_/X _18393_/A _18391_/X VGND VGND VPWR VPWR _18392_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17338_/A _17317_/C _17288_/X _17340_/B VGND VGND VPWR VPWR _17343_/X sky130_fd_sc_hd__a211o_4
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ _23971_/Q _14555_/B VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__and2_4
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11765_/Y _11760_/X _11766_/X _11760_/X VGND VGND VPWR VPWR _11767_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21151__A1 _13526_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13506_/A VGND VGND VPWR VPWR _13516_/A sky130_fd_sc_hd__inv_2
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17274_/A _17271_/A VGND VGND VPWR VPWR _17274_/X sky130_fd_sc_hd__or2_4
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _14483_/Y _14485_/X _14420_/X _14485_/X VGND VGND VPWR VPWR _25126_/D sky130_fd_sc_hd__a2bb2o_4
X_11698_ _13740_/B VGND VGND VPWR VPWR _13690_/B sky130_fd_sc_hd__inv_2
XFILLER_146_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19013_ _19020_/A VGND VGND VPWR VPWR _19013_/X sky130_fd_sc_hd__buf_2
X_16225_ _16224_/Y _16222_/X _15965_/X _16222_/X VGND VGND VPWR VPWR _16225_/X sky130_fd_sc_hd__a2bb2o_4
X_13437_ _13469_/A _13435_/X _13437_/C VGND VGND VPWR VPWR _13438_/C sky130_fd_sc_hd__and3_4
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17728__A2_N _21675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16156_ _24694_/Q VGND VGND VPWR VPWR _16156_/Y sky130_fd_sc_hd__inv_2
X_13368_ _13243_/X _13368_/B VGND VGND VPWR VPWR _13368_/X sky130_fd_sc_hd__or2_4
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15107_ _24989_/Q VGND VGND VPWR VPWR _15411_/A sky130_fd_sc_hd__inv_2
X_12319_ _25361_/Q _12317_/Y _12306_/A _12318_/Y VGND VGND VPWR VPWR _12322_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16087_ _11730_/Y _21299_/A _15933_/X _21071_/A _16086_/X VGND VGND VPWR VPWR _24720_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_181_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21984__B _21983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13299_ _13178_/A _13299_/B VGND VGND VPWR VPWR _13299_/X sky130_fd_sc_hd__or2_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15038_ _25017_/Q _15036_/Y _25019_/Q _15037_/Y VGND VGND VPWR VPWR _15042_/C sky130_fd_sc_hd__a2bb2o_4
X_19915_ _19914_/Y _19910_/X _19639_/X _19910_/X VGND VGND VPWR VPWR _19915_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18607__B1 _16550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25141__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20414__B1 _20243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19846_ _23609_/Q VGND VGND VPWR VPWR _21894_/B sky130_fd_sc_hd__inv_2
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16989_ _16982_/X _16984_/X _16989_/C _16988_/X VGND VGND VPWR VPWR _16989_/X sky130_fd_sc_hd__or4_4
X_19777_ _13371_/B VGND VGND VPWR VPWR _19777_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12399__A _12391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19296__A2_N _19293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_252_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _23980_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15841__B1 _15632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14911__A1_N _25023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18728_ _18739_/A _18726_/X _18728_/C VGND VGND VPWR VPWR _24158_/D sky130_fd_sc_hd__and3_4
XFILLER_25_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21505__A _21668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18659_ _18659_/A _18659_/B _18659_/C _18659_/D VGND VGND VPWR VPWR _18659_/X sky130_fd_sc_hd__or4_4
XFILLER_92_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15503__A _15503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21670_ _21482_/A _21670_/B _21669_/X VGND VGND VPWR VPWR _21670_/X sky130_fd_sc_hd__and3_4
XFILLER_197_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20621_ _13976_/A _20621_/B _15438_/C VGND VGND VPWR VPWR _23978_/D sky130_fd_sc_hd__and3_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23340_ _22810_/A _23339_/Y VGND VGND VPWR VPWR _23340_/Y sky130_fd_sc_hd__nor2_4
X_20552_ _20552_/A _18893_/A VGND VGND VPWR VPWR _20552_/X sky130_fd_sc_hd__and2_4
XFILLER_193_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23271_ _16657_/Y _22842_/X _15574_/Y _22845_/X VGND VGND VPWR VPWR _23271_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20483_ _20503_/B VGND VGND VPWR VPWR _20682_/B sky130_fd_sc_hd__buf_2
XANTENNA__16334__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22222_ _21262_/A _22214_/X _22221_/X VGND VGND VPWR VPWR _22222_/X sky130_fd_sc_hd__and3_4
X_25010_ _25011_/CLK _25010_/D HRESETn VGND VGND VPWR VPWR _25010_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22642__A1 _21058_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18846__B1 _16524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24343__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22642__B2 _22565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22153_ _22947_/A VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__buf_2
X_21104_ _24617_/Q _21104_/B VGND VGND VPWR VPWR _21104_/X sky130_fd_sc_hd__or2_4
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22084_ _22079_/X _22083_/X _14686_/X VGND VGND VPWR VPWR _22084_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22071__A _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14883__A1 _14877_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_62_0_HCLK clkbuf_5_31_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _21035_/A _21034_/X VGND VGND VPWR VPWR _21060_/B sky130_fd_sc_hd__or2_4
XFILLER_247_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16085__B1 _15489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24856__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22158__B1 _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15832__B1 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19023__B1 _18908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22986_ _22986_/A VGND VGND VPWR VPWR _22986_/X sky130_fd_sc_hd__buf_2
XFILLER_228_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24725_ _24726_/CLK _16077_/X HRESETn VGND VGND VPWR VPWR _24725_/Q sky130_fd_sc_hd__dfrtp_4
X_21937_ _21941_/A _21937_/B VGND VGND VPWR VPWR _21939_/B sky130_fd_sc_hd__or2_4
XFILLER_215_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12131__A1_N _12175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12670_ _12628_/X _12647_/D _12588_/Y VGND VGND VPWR VPWR _12671_/C sky130_fd_sc_hd__o21a_4
X_24656_ _24169_/CLK _24656_/D HRESETn VGND VGND VPWR VPWR _16268_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_230_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21868_ _17250_/A _21868_/B VGND VGND VPWR VPWR _21868_/X sky130_fd_sc_hd__or2_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _24295_/CLK _19852_/X VGND VGND VPWR VPWR _19850_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_169_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20822_/B _13145_/X _20818_/X VGND VGND VPWR VPWR _20819_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _14730_/C _22062_/A VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__and2_4
X_24587_ _24989_/CLK _24587_/D HRESETn VGND VGND VPWR VPWR _15124_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17050__D _17050_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18724__A _18710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _25173_/Q _14369_/A _14335_/X VGND VGND VPWR VPWR _14340_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23538_ _23560_/CLK _20045_/X VGND VGND VPWR VPWR _20043_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15899__B1 _22726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271_ _14270_/Y _14268_/X _13846_/X _14268_/X VGND VGND VPWR VPWR _14271_/X sky130_fd_sc_hd__a2bb2o_4
X_23469_ _23493_/CLK _20231_/X VGND VGND VPWR VPWR _23469_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16010_ _16010_/A VGND VGND VPWR VPWR _16010_/Y sky130_fd_sc_hd__inv_2
X_13222_ _13320_/A VGND VGND VPWR VPWR _13222_/X sky130_fd_sc_hd__buf_2
X_25208_ _25253_/CLK _25208_/D HRESETn VGND VGND VPWR VPWR _14223_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22633__B2 _21322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ _13211_/A VGND VGND VPWR VPWR _13153_/X sky130_fd_sc_hd__buf_2
X_25139_ _25223_/CLK _14454_/X HRESETn VGND VGND VPWR VPWR _25139_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15115__A2 _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12104_ _21031_/A VGND VGND VPWR VPWR _17448_/A sky130_fd_sc_hd__inv_2
X_13084_ _13006_/A _13084_/B VGND VGND VPWR VPWR _13085_/C sky130_fd_sc_hd__or2_4
X_17961_ _17957_/X _17960_/X _18027_/A VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__o21a_4
XFILLER_239_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24128__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _12035_/A _12027_/X _12035_/C _12034_/X VGND VGND VPWR VPWR _14299_/B sky130_fd_sc_hd__or4_4
X_16912_ _16175_/Y _21066_/A _16175_/Y _21066_/A VGND VGND VPWR VPWR _16912_/X sky130_fd_sc_hd__a2bb2o_4
X_19700_ _19696_/Y _19699_/X _19677_/X _19699_/X VGND VGND VPWR VPWR _19700_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17892_ _17881_/A _17888_/X _17892_/C VGND VGND VPWR VPWR _17892_/X sky130_fd_sc_hd__and3_4
XFILLER_78_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24597__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16843_ _16843_/A VGND VGND VPWR VPWR _16843_/Y sky130_fd_sc_hd__inv_2
X_19631_ _23682_/Q VGND VGND VPWR VPWR _19631_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13753__D _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15823__B1 _11797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19562_ _23704_/Q VGND VGND VPWR VPWR _19562_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19014__B1 _19012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16774_ _16772_/Y _16768_/X _15754_/X _16773_/X VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__a2bb2o_4
X_13986_ _25238_/Q VGND VGND VPWR VPWR _14027_/A sky130_fd_sc_hd__buf_2
XFILLER_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18513_ _18828_/B _18513_/B _18512_/X VGND VGND VPWR VPWR _18514_/A sky130_fd_sc_hd__or3_4
X_15725_ _15725_/A VGND VGND VPWR VPWR _15772_/A sky130_fd_sc_hd__inv_2
X_12937_ _12927_/A _12935_/X _12936_/X VGND VGND VPWR VPWR _25388_/D sky130_fd_sc_hd__and3_4
X_19493_ _19493_/A VGND VGND VPWR VPWR _21825_/B sky130_fd_sc_hd__inv_2
XFILLER_206_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16419__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_82_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24799_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11851__A _11851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18444_ _16219_/Y _24185_/Q _22557_/A _18479_/D VGND VGND VPWR VPWR _18451_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15656_ _13818_/A VGND VGND VPWR VPWR _15656_/X sky130_fd_sc_hd__buf_2
XFILLER_222_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21044__B _21069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12868_ _25404_/Q _12868_/B VGND VGND VPWR VPWR _12868_/X sky130_fd_sc_hd__or2_4
XPHY_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14607_/A _14574_/B VGND VGND VPWR VPWR _14607_/Y sky130_fd_sc_hd__nand2_4
X_11819_ _11816_/Y _11814_/X _11818_/X _11814_/X VGND VGND VPWR VPWR _11819_/X sky130_fd_sc_hd__a2bb2o_4
X_18375_ _18374_/Y _18362_/Y _18372_/A _18361_/X VGND VGND VPWR VPWR _18375_/X sky130_fd_sc_hd__o22a_4
X_15587_ _15586_/Y _15584_/X _11776_/X _15584_/X VGND VGND VPWR VPWR _15587_/X sky130_fd_sc_hd__a2bb2o_4
X_12799_ _12799_/A _12799_/B _12799_/C _12798_/X VGND VGND VPWR VPWR _12799_/X sky130_fd_sc_hd__or4_4
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17326_ _17331_/A _17330_/A _17262_/Y _17326_/D VGND VGND VPWR VPWR _17332_/B sky130_fd_sc_hd__or4_4
XANTENNA__17879__A1 _16920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14538_ _14530_/X _14537_/X _25121_/Q _14515_/Y VGND VGND VPWR VPWR _25109_/D sky130_fd_sc_hd__o22a_4
XFILLER_175_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_202_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22156__A _21300_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17257_ _17348_/A VGND VGND VPWR VPWR _17257_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14469_ _14467_/Y _14463_/X _14427_/X _14468_/X VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16208_ _16207_/Y _16203_/X _15952_/X _16203_/X VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__a2bb2o_4
X_17188_ _24638_/Q _17322_/A _24644_/Q _17294_/A VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16139_ _16138_/Y _16136_/X _11809_/X _16136_/X VGND VGND VPWR VPWR _16139_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15993__A _11861_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20938__A1 _16671_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16067__B1 _16066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19829_ _19816_/A VGND VGND VPWR VPWR _19829_/X sky130_fd_sc_hd__buf_2
XFILLER_217_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15814__B1 _24850_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19005__B1 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22840_ _12819_/Y _21456_/X _17832_/A _22839_/X VGND VGND VPWR VPWR _22840_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21880__D _21879_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22771_ _21890_/X VGND VGND VPWR VPWR _22771_/X sky130_fd_sc_hd__buf_2
XANTENNA__12857__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24510_ _24509_/CLK _16665_/X HRESETn VGND VGND VPWR VPWR _16664_/A sky130_fd_sc_hd__dfrtp_4
X_21722_ _12273_/X _21542_/A _24266_/Q _21440_/X VGND VGND VPWR VPWR _21724_/A sky130_fd_sc_hd__a2bb2o_4
X_25490_ _25491_/CLK _12086_/X HRESETn VGND VGND VPWR VPWR _12085_/A sky130_fd_sc_hd__dfrtp_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23104__A2 _23095_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12575__A2_N _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _13826_/X VGND VGND VPWR VPWR _22549_/B sky130_fd_sc_hd__buf_2
X_24441_ _24437_/CLK _16824_/X HRESETn VGND VGND VPWR VPWR _14980_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20604_ _23961_/Q _18888_/B _18890_/A VGND VGND VPWR VPWR _20604_/Y sky130_fd_sc_hd__a21oi_4
X_21584_ _21583_/X VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__buf_2
X_24372_ _24372_/CLK _17299_/Y HRESETn VGND VGND VPWR VPWR _17245_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20535_ _20535_/A _20503_/X _20510_/X _20527_/A VGND VGND VPWR VPWR _20535_/X sky130_fd_sc_hd__or4_4
X_23323_ _21881_/X _23322_/X _22484_/X _24891_/Q _21085_/A VGND VGND VPWR VPWR _23324_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_138_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20466_ _20438_/A _20464_/X _20460_/A _20465_/X VGND VGND VPWR VPWR _20466_/Y sky130_fd_sc_hd__a22oi_4
X_23254_ _24613_/Q _23313_/B VGND VGND VPWR VPWR _23254_/X sky130_fd_sc_hd__or2_4
X_22205_ _22171_/X _22205_/B _22205_/C _22204_/X VGND VGND VPWR VPWR _22205_/X sky130_fd_sc_hd__or4_4
X_23185_ _16482_/A _23184_/X _23148_/X VGND VGND VPWR VPWR _23185_/X sky130_fd_sc_hd__o21a_4
XFILLER_145_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20397_ _23406_/Q VGND VGND VPWR VPWR _21682_/B sky130_fd_sc_hd__inv_2
XFILLER_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22513__B _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22136_ _21350_/Y _22119_/X _22123_/Y _22128_/Y _22135_/X VGND VGND VPWR VPWR _22136_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_160_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22067_ _25265_/Q _22524_/B _13792_/A _22066_/Y VGND VGND VPWR VPWR _22067_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19244__B1 _19220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17326__C _17262_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24690__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21018_ _21018_/A _21018_/B VGND VGND VPWR VPWR _21018_/Y sky130_fd_sc_hd__nor2_4
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15805__B1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13840_ _13840_/A VGND VGND VPWR VPWR _13840_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23343__A2 _22485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13771_ _13770_/X VGND VGND VPWR VPWR _13771_/X sky130_fd_sc_hd__buf_2
XFILLER_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22969_ _14978_/A _22851_/X _22108_/X _22968_/X VGND VGND VPWR VPWR _22969_/X sky130_fd_sc_hd__a211o_4
XFILLER_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17558__B1 _11853_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22551__B1 _21968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15510_ _11736_/B VGND VGND VPWR VPWR _15510_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_69_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12722_ _12728_/A _12722_/B _12722_/C VGND VGND VPWR VPWR _12722_/X sky130_fd_sc_hd__and3_4
X_24708_ _24712_/CLK _24708_/D HRESETn VGND VGND VPWR VPWR _24708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16490_ _24575_/Q VGND VGND VPWR VPWR _16490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16230__B1 _15970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15441_ _15440_/X VGND VGND VPWR VPWR _15441_/X sky130_fd_sc_hd__buf_2
X_12653_ _25433_/Q _12657_/B VGND VGND VPWR VPWR _12655_/B sky130_fd_sc_hd__or2_4
X_24639_ _24639_/CLK _16318_/X HRESETn VGND VGND VPWR VPWR _16317_/A sky130_fd_sc_hd__dfrtp_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21106__A1 _24650_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ _18060_/A _23775_/Q VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__or2_4
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _15305_/A _15377_/B _15348_/X VGND VGND VPWR VPWR _15372_/Y sky130_fd_sc_hd__a21oi_4
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12619_/B _12568_/A _25427_/Q _12535_/Y VGND VGND VPWR VPWR _12584_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _16996_/Y _17118_/A _17042_/B _17120_/B VGND VGND VPWR VPWR _17117_/B sky130_fd_sc_hd__or4_4
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _14315_/X _14322_/X _13490_/A _14320_/X VGND VGND VPWR VPWR _14323_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13598__A _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18091_ _18126_/A _23881_/Q VGND VGND VPWR VPWR _18092_/C sky130_fd_sc_hd__or2_4
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17042_ _16981_/Y _17042_/B _17042_/C _17042_/D VGND VGND VPWR VPWR _17042_/X sky130_fd_sc_hd__or4_4
X_14254_ _14254_/A _14254_/B VGND VGND VPWR VPWR _14255_/B sky130_fd_sc_hd__or2_4
XANTENNA__22606__A1 _22563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22606__B2 _22565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13205_ _13267_/A VGND VGND VPWR VPWR _13207_/A sky130_fd_sc_hd__inv_2
X_14185_ _14185_/A VGND VGND VPWR VPWR _14185_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24778__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _13136_/A _13136_/B VGND VGND VPWR VPWR _13137_/B sky130_fd_sc_hd__or2_4
X_18993_ _18990_/Y _18986_/X _18991_/X _18992_/X VGND VGND VPWR VPWR _18993_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24707__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11846__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13067_ _13063_/B _13066_/X VGND VGND VPWR VPWR _13068_/B sky130_fd_sc_hd__or2_4
X_17944_ _17944_/A _19001_/A VGND VGND VPWR VPWR _17945_/C sky130_fd_sc_hd__or2_4
XFILLER_239_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12018_ _24106_/Q _12001_/X _12017_/Y VGND VGND VPWR VPWR _12019_/A sky130_fd_sc_hd__o21a_4
X_17875_ _17875_/A VGND VGND VPWR VPWR _17875_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19614_ _19614_/A VGND VGND VPWR VPWR _19614_/Y sky130_fd_sc_hd__inv_2
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16826_ _14913_/Y _16825_/X HWDATA[21] _16825_/X VGND VGND VPWR VPWR _16826_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23254__B _23313_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21055__A _21046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16757_ _16756_/Y _16752_/X _16407_/X _16752_/X VGND VGND VPWR VPWR _24473_/D sky130_fd_sc_hd__a2bb2o_4
X_19545_ _23709_/Q VGND VGND VPWR VPWR _21192_/B sky130_fd_sc_hd__inv_2
X_13969_ _13969_/A VGND VGND VPWR VPWR _13969_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15708_ _24892_/Q _15707_/X _15699_/X VGND VGND VPWR VPWR _15708_/X sky130_fd_sc_hd__o21a_4
X_16688_ _16687_/Y _16685_/X _16419_/X _16685_/X VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__a2bb2o_4
X_19476_ _19475_/Y _19473_/X _19454_/X _19473_/X VGND VGND VPWR VPWR _19476_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15639_ _15638_/Y _15635_/X _15480_/X _15635_/X VGND VGND VPWR VPWR _24902_/D sky130_fd_sc_hd__a2bb2o_4
X_18427_ _24181_/Q VGND VGND VPWR VPWR _18540_/A sky130_fd_sc_hd__inv_2
XFILLER_221_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18358_ _18357_/Y _17487_/Y _18357_/A _17492_/X VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__o22a_4
X_17309_ _17300_/X VGND VGND VPWR VPWR _17313_/B sky130_fd_sc_hd__inv_2
XFILLER_147_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18289_ _18289_/A _18288_/X _18289_/C VGND VGND VPWR VPWR _18289_/X sky130_fd_sc_hd__or3_4
XFILLER_163_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20320_ _21200_/B _20315_/X _20034_/X _20302_/Y VGND VGND VPWR VPWR _20320_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20251_ _18178_/B VGND VGND VPWR VPWR _20251_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23270__B2 _22298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20182_ _20181_/Y _20177_/X _20115_/X _20177_/X VGND VGND VPWR VPWR _23488_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24990_ _24966_/CLK _24990_/D HRESETn VGND VGND VPWR VPWR _24990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23941_ _25106_/CLK _23941_/D HRESETn VGND VGND VPWR VPWR _23941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23872_ _23871_/CLK _19088_/X VGND VGND VPWR VPWR _13346_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22823_ _22944_/A _22823_/B _22822_/X VGND VGND VPWR VPWR _22824_/D sky130_fd_sc_hd__and3_4
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21336__A1 _24452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25542_ _25539_/CLK _25542_/D HRESETn VGND VGND VPWR VPWR _25542_/Q sky130_fd_sc_hd__dfrtp_4
X_22754_ _22754_/A _22754_/B _22754_/C VGND VGND VPWR VPWR _22754_/X sky130_fd_sc_hd__and3_4
XFILLER_197_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21705_ _18278_/X _21703_/X _21520_/X _21704_/Y VGND VGND VPWR VPWR _21706_/A sky130_fd_sc_hd__a211o_4
X_25473_ _24112_/CLK _12173_/X HRESETn VGND VGND VPWR VPWR _18377_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22685_ _16599_/Y _23027_/B _21591_/X _22684_/X VGND VGND VPWR VPWR _22685_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24424_ _24425_/CLK _16855_/X HRESETn VGND VGND VPWR VPWR _14954_/A sky130_fd_sc_hd__dfrtp_4
X_21636_ _22090_/A _19937_/Y VGND VGND VPWR VPWR _21636_/X sky130_fd_sc_hd__or2_4
XFILLER_185_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11815__A1_N _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24355_ _25494_/CLK _17371_/X HRESETn VGND VGND VPWR VPWR _24355_/Q sky130_fd_sc_hd__dfrtp_4
X_21567_ _21567_/A _21733_/B VGND VGND VPWR VPWR _21567_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23306_ _23136_/X _23306_/B VGND VGND VPWR VPWR _23306_/Y sky130_fd_sc_hd__nor2_4
XFILLER_181_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20518_ _20518_/A _20684_/A VGND VGND VPWR VPWR _20518_/X sky130_fd_sc_hd__and2_4
X_21498_ _21808_/A _21498_/B _21497_/X VGND VGND VPWR VPWR _21498_/X sky130_fd_sc_hd__and3_4
X_24286_ _24272_/CLK _24286_/D HRESETn VGND VGND VPWR VPWR _17751_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20449_ _20449_/A VGND VGND VPWR VPWR _20451_/A sky130_fd_sc_hd__inv_2
X_23237_ _23237_/A _23296_/B VGND VGND VPWR VPWR _23237_/X sky130_fd_sc_hd__or2_4
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16522__A _16522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16279__B1 _15489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24871__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20075__B2 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23168_ _22204_/A VGND VGND VPWR VPWR _23168_/X sky130_fd_sc_hd__buf_2
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24800__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ _22119_/A _22114_/Y _22119_/C _22118_/X VGND VGND VPWR VPWR _22119_/X sky130_fd_sc_hd__or4_4
X_15990_ _15945_/Y VGND VGND VPWR VPWR _15990_/X sky130_fd_sc_hd__buf_2
X_23099_ _23099_/A VGND VGND VPWR VPWR _23099_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14941_ _15270_/A VGND VGND VPWR VPWR _15072_/A sky130_fd_sc_hd__inv_2
XFILLER_248_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21575__B2 _16731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17660_ _17644_/A _17635_/X _17611_/X _17658_/B VGND VGND VPWR VPWR _17661_/A sky130_fd_sc_hd__a211o_4
X_14872_ _14852_/A _14871_/Y _14822_/C _14852_/A VGND VGND VPWR VPWR _25050_/D sky130_fd_sc_hd__a2bb2o_4
X_16611_ _16608_/Y _16604_/X _16609_/X _16610_/X VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__a2bb2o_4
X_13823_ _14415_/A _14462_/A VGND VGND VPWR VPWR _17422_/A sky130_fd_sc_hd__or2_4
X_17591_ _17621_/D _17590_/X VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__or2_4
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16542_ _16542_/A VGND VGND VPWR VPWR _16542_/Y sky130_fd_sc_hd__inv_2
X_19330_ _19330_/A VGND VGND VPWR VPWR _19330_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13754_ _13753_/X VGND VGND VPWR VPWR _13754_/X sky130_fd_sc_hd__buf_2
XANTENNA__21878__A2 _22299_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ _25419_/Q _12705_/B VGND VGND VPWR VPWR _12705_/X sky130_fd_sc_hd__or2_4
X_19261_ _23811_/Q VGND VGND VPWR VPWR _19261_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16473_ _16472_/Y _16470_/X _16294_/X _16470_/X VGND VGND VPWR VPWR _24582_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13685_ _25301_/Q VGND VGND VPWR VPWR _13685_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18212_ _18051_/A _18208_/X _18212_/C VGND VGND VPWR VPWR _18220_/B sky130_fd_sc_hd__or3_4
X_15424_ _15424_/A _15424_/B VGND VGND VPWR VPWR _15424_/X sky130_fd_sc_hd__or2_4
XFILLER_231_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22418__B _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12636_ _12636_/A _12634_/X _12635_/X VGND VGND VPWR VPWR _25437_/D sky130_fd_sc_hd__and3_4
X_19192_ _19188_/Y _19191_/X _19169_/X _19191_/X VGND VGND VPWR VPWR _19192_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_156_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24196_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _18036_/A _18143_/B VGND VGND VPWR VPWR _18143_/X sky130_fd_sc_hd__or2_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _15355_/A _15346_/X _15355_/C VGND VGND VPWR VPWR _25004_/D sky130_fd_sc_hd__and3_4
XFILLER_8_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12567_ _12567_/A _12540_/X _12553_/X _12566_/X VGND VGND VPWR VPWR _12609_/A sky130_fd_sc_hd__or4_4
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _14300_/A _14305_/X _13649_/X VGND VGND VPWR VPWR _14306_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_144_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18074_ _18036_/A _18074_/B VGND VGND VPWR VPWR _18074_/X sky130_fd_sc_hd__or2_4
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15286_ _15292_/A _15256_/X VGND VGND VPWR VPWR _15293_/B sky130_fd_sc_hd__or2_4
X_12498_ _12218_/Y _12501_/B _12403_/X VGND VGND VPWR VPWR _12498_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_144_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17025_ _17021_/X _17022_/X _17025_/C _17024_/X VGND VGND VPWR VPWR _17025_/X sky130_fd_sc_hd__or4_4
X_14237_ _20672_/A VGND VGND VPWR VPWR _14237_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16432__A _16432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20066__B2 _20065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ _14108_/C _14122_/X _14108_/C _14122_/X VGND VGND VPWR VPWR _14169_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ _13117_/Y _13118_/X _13121_/C VGND VGND VPWR VPWR _13119_/X sky130_fd_sc_hd__and3_4
XANTENNA__19208__B1 _19139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19743__A _19742_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _20549_/B _14556_/B _14078_/X _13994_/B _14093_/X VGND VGND VPWR VPWR _25233_/D
+ sky130_fd_sc_hd__a32o_4
X_18976_ _18973_/Y _18974_/X _18975_/X _18974_/X VGND VGND VPWR VPWR _23911_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16690__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17927_ _17921_/Y _13550_/X _17924_/Y _24258_/Q _17926_/X VGND VGND VPWR VPWR _17927_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17263__A _17331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17858_ _17759_/X _17858_/B VGND VGND VPWR VPWR _17858_/X sky130_fd_sc_hd__or2_4
XFILLER_226_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16809_ _16808_/Y _16806_/X _15723_/X _16806_/X VGND VGND VPWR VPWR _16809_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21318__A1 _21307_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17789_ _17748_/X _17789_/B _17789_/C VGND VGND VPWR VPWR _17789_/X sky130_fd_sc_hd__and3_4
XFILLER_19_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19528_ _19527_/X VGND VGND VPWR VPWR _19528_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_52_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19459_ _14665_/Y _13634_/X _19028_/C VGND VGND VPWR VPWR _19460_/A sky130_fd_sc_hd__or3_4
XFILLER_179_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14756__B1 _14725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _12113_/Y _12081_/B _12023_/Y _13484_/D VGND VGND VPWR VPWR _22470_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21232__B _21877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21421_ _14723_/A _21413_/X _21420_/X VGND VGND VPWR VPWR _21421_/X sky130_fd_sc_hd__or3_4
XANTENNA__19695__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21352_ _21352_/A _22190_/B VGND VGND VPWR VPWR _21361_/A sky130_fd_sc_hd__and2_4
X_24140_ _25212_/CLK _18806_/X HRESETn VGND VGND VPWR VPWR _24140_/Q sky130_fd_sc_hd__dfrtp_4
X_20303_ _20302_/Y VGND VGND VPWR VPWR _20303_/X sky130_fd_sc_hd__buf_2
XANTENNA__24629__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21283_ _21384_/B _21281_/X _25276_/Q _21282_/X VGND VGND VPWR VPWR _21283_/X sky130_fd_sc_hd__o22a_4
X_24071_ _24073_/CLK _24071_/D HRESETn VGND VGND VPWR VPWR _20944_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__19447__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20234_ _20233_/X VGND VGND VPWR VPWR _20234_/Y sky130_fd_sc_hd__inv_2
X_23022_ _16219_/A _22827_/B VGND VGND VPWR VPWR _23025_/B sky130_fd_sc_hd__or2_4
XFILLER_116_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20165_ _23494_/Q VGND VGND VPWR VPWR _20165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19653__A _19652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15487__A1_N _14877_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16681__B1 _16412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20096_ _20095_/Y _20093_/X _19832_/X _20093_/X VGND VGND VPWR VPWR _20096_/X sky130_fd_sc_hd__a2bb2o_4
X_24973_ _24966_/CLK _15457_/X HRESETn VGND VGND VPWR VPWR _13950_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21557__A1 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23924_ _25491_/CLK _18941_/X VGND VGND VPWR VPWR _23924_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18422__A1 _16201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16433__B1 _16248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23855_ _23871_/CLK _19135_/X VGND VGND VPWR VPWR _23855_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22806_ _22801_/X _22803_/X _22804_/X _22805_/X VGND VGND VPWR VPWR _22807_/B sky130_fd_sc_hd__o22a_4
XFILLER_44_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23786_ _24252_/CLK _23786_/D VGND VGND VPWR VPWR _19330_/A sky130_fd_sc_hd__dfxtp_4
X_20998_ _20998_/A VGND VGND VPWR VPWR _21000_/B sky130_fd_sc_hd__inv_2
XFILLER_213_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25525_ _24386_/CLK _25525_/D HRESETn VGND VGND VPWR VPWR _25525_/Q sky130_fd_sc_hd__dfrtp_4
X_22737_ _22737_/A _22737_/B _22729_/X _22736_/Y VGND VGND VPWR VPWR HRDATA[14] sky130_fd_sc_hd__or4_4
XFILLER_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25070__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13470_ _13332_/X _13466_/X _13470_/C VGND VGND VPWR VPWR _13471_/C sky130_fd_sc_hd__or3_4
X_25456_ _25456_/CLK _12455_/X HRESETn VGND VGND VPWR VPWR _12208_/A sky130_fd_sc_hd__dfrtp_4
X_22668_ _21090_/A VGND VGND VPWR VPWR _22669_/B sky130_fd_sc_hd__buf_2
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_229_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24138_/CLK sky130_fd_sc_hd__clkbuf_1
X_12421_ _12421_/A _12415_/Y _12421_/C VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__or3_4
X_24407_ _24407_/CLK _24407_/D HRESETn VGND VGND VPWR VPWR _16990_/A sky130_fd_sc_hd__dfrtp_4
X_21619_ _22235_/A VGND VGND VPWR VPWR _21646_/A sky130_fd_sc_hd__buf_2
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25387_ _25402_/CLK _25387_/D HRESETn VGND VGND VPWR VPWR _22724_/A sky130_fd_sc_hd__dfrtp_4
X_22599_ _22528_/X _22596_/X _22431_/X _22598_/X VGND VGND VPWR VPWR _22599_/X sky130_fd_sc_hd__o22a_4
X_15140_ _15139_/Y _16427_/A _15139_/Y _16427_/A VGND VGND VPWR VPWR _15141_/D sky130_fd_sc_hd__a2bb2o_4
X_12352_ _25357_/Q _12350_/Y _12351_/Y _24830_/Q VGND VGND VPWR VPWR _12360_/A sky130_fd_sc_hd__a2bb2o_4
X_24338_ _25200_/CLK _17428_/X HRESETn VGND VGND VPWR VPWR _20675_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_193_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15071_ _14990_/A _15290_/A _15292_/A VGND VGND VPWR VPWR _15071_/X sky130_fd_sc_hd__or3_4
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12283_ _12282_/X VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__buf_2
X_24269_ _24715_/CLK _24269_/D HRESETn VGND VGND VPWR VPWR _22199_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16252__A _16252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14022_ _14022_/A _14022_/B VGND VGND VPWR VPWR _14556_/A sky130_fd_sc_hd__nor2_4
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21796__B2 _21656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18830_ pwm_S7 VGND VGND VPWR VPWR _18830_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15973_ _12237_/Y _15968_/X _15972_/X _15968_/X VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__a2bb2o_4
X_18761_ _18698_/C _18766_/B _18714_/X VGND VGND VPWR VPWR _18761_/Y sky130_fd_sc_hd__a21oi_4
X_14924_ _14924_/A VGND VGND VPWR VPWR _15016_/A sky130_fd_sc_hd__inv_2
X_17712_ _17712_/A VGND VGND VPWR VPWR _17898_/B sky130_fd_sc_hd__inv_2
XFILLER_48_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18692_ _18782_/A VGND VGND VPWR VPWR _18699_/A sky130_fd_sc_hd__inv_2
XANTENNA__16424__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20220__B2 _20219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14855_ _25055_/Q _14824_/X _25055_/Q _14824_/X VGND VGND VPWR VPWR _14856_/A sky130_fd_sc_hd__a2bb2o_4
X_17643_ _17642_/X VGND VGND VPWR VPWR _24316_/D sky130_fd_sc_hd__inv_2
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15778__A2 _15774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13806_ _14400_/A VGND VGND VPWR VPWR _13806_/X sky130_fd_sc_hd__buf_2
X_17574_ _24312_/Q VGND VGND VPWR VPWR _17646_/C sky130_fd_sc_hd__inv_2
XFILLER_205_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14786_ _14783_/A _14785_/A _14772_/A _14781_/A VGND VGND VPWR VPWR _14787_/A sky130_fd_sc_hd__a211o_4
X_11998_ _25500_/Q VGND VGND VPWR VPWR _11998_/Y sky130_fd_sc_hd__inv_2
X_16525_ _16533_/A VGND VGND VPWR VPWR _16525_/X sky130_fd_sc_hd__buf_2
X_19313_ _23792_/Q VGND VGND VPWR VPWR _19313_/Y sky130_fd_sc_hd__inv_2
X_13737_ _13692_/X _13736_/Y _13730_/X _13722_/X _11678_/A VGND VGND VPWR VPWR _25289_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_39_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16427__A _16427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22148__B _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21720__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16456_ _24584_/Q VGND VGND VPWR VPWR _18515_/A sky130_fd_sc_hd__inv_2
X_19244_ _19243_/Y _19241_/X _19220_/X _19241_/X VGND VGND VPWR VPWR _23817_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13668_ _20865_/A _20865_/B _24056_/Q _24055_/Q VGND VGND VPWR VPWR _13668_/X sky130_fd_sc_hd__or4_4
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15407_ _15407_/A _15407_/B VGND VGND VPWR VPWR _15408_/C sky130_fd_sc_hd__nand2_4
X_12619_ _12619_/A _12619_/B _12618_/X VGND VGND VPWR VPWR _12620_/C sky130_fd_sc_hd__or3_4
X_19175_ _19173_/Y _19168_/X _19151_/X _19174_/X VGND VGND VPWR VPWR _19175_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16387_ _16387_/A VGND VGND VPWR VPWR _16387_/Y sky130_fd_sc_hd__inv_2
X_13599_ _13551_/X _13599_/B VGND VGND VPWR VPWR _14629_/B sky130_fd_sc_hd__and2_4
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12359__A2_N _24839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24793__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18126_ _18126_/A _19065_/A VGND VGND VPWR VPWR _18127_/C sky130_fd_sc_hd__or2_4
XFILLER_191_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15338_ _15340_/B VGND VGND VPWR VPWR _15343_/B sky130_fd_sc_hd__inv_2
XANTENNA__20287__B2 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24722__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _18130_/A _18055_/X _18057_/C VGND VGND VPWR VPWR _18057_/X sky130_fd_sc_hd__and3_4
XANTENNA__13786__A _13786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _15271_/B VGND VGND VPWR VPWR _15270_/B sky130_fd_sc_hd__inv_2
XFILLER_172_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ _16051_/Y _17045_/A _16051_/Y _17045_/A VGND VGND VPWR VPWR _17008_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19473__A _19460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16663__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18959_ _18959_/A _18959_/B _18938_/A _18938_/B VGND VGND VPWR VPWR _18959_/X sky130_fd_sc_hd__or4_4
XFILLER_101_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22197__D1 _22196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21970_ _25264_/Q _13824_/X VGND VGND VPWR VPWR _21970_/X sky130_fd_sc_hd__or2_4
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20921_ _16682_/Y _20854_/A _20863_/X _20920_/Y VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23640_ _23631_/CLK _23640_/D VGND VGND VPWR VPWR _13369_/B sky130_fd_sc_hd__dfxtp_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _16718_/Y _20833_/X _20842_/X _20851_/Y VGND VGND VPWR VPWR _20852_/X sky130_fd_sc_hd__o22a_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21243__A _21267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23571_ _23529_/CLK _23571_/D VGND VGND VPWR VPWR _19948_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20783_ _20782_/X VGND VGND VPWR VPWR _20783_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12865__A _12638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25310_ _23631_/CLK _13540_/X HRESETn VGND VGND VPWR VPWR SCLK_S2 sky130_fd_sc_hd__dfstp_4
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22522_ _22522_/A VGND VGND VPWR VPWR _22536_/B sky130_fd_sc_hd__inv_2
XFILLER_222_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25241_ _25246_/CLK _25241_/D HRESETn VGND VGND VPWR VPWR _13999_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22453_ _22306_/A VGND VGND VPWR VPWR _22453_/X sky130_fd_sc_hd__buf_2
XFILLER_195_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21404_ _14700_/X _21402_/X _21403_/X VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__and3_4
X_25172_ _25168_/CLK _14343_/X HRESETn VGND VGND VPWR VPWR _25172_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22384_ _22380_/X _22383_/X _14686_/X VGND VGND VPWR VPWR _22384_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24123_ _25106_/CLK _18900_/X HRESETn VGND VGND VPWR VPWR _21000_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_59_0_HCLK clkbuf_8_58_0_HCLK/A VGND VGND VPWR VPWR _25281_/CLK sky130_fd_sc_hd__clkbuf_1
X_21335_ _21334_/Y VGND VGND VPWR VPWR _21335_/X sky130_fd_sc_hd__buf_2
XANTENNA__23216__B2 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16072__A _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24054_ _24493_/CLK _24054_/D HRESETn VGND VGND VPWR VPWR _20865_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21266_ _21273_/A _19878_/Y VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__or2_4
XANTENNA__22802__A _22694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22975__B1 _11789_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23005_ _23072_/A _23005_/B VGND VGND VPWR VPWR _23005_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24959__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20217_ _20216_/Y _20214_/X _16870_/X _20214_/X VGND VGND VPWR VPWR _20217_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19383__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21197_ _21193_/X _21196_/X _24219_/Q VGND VGND VPWR VPWR _21197_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15457__A1 _14289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20148_ _23500_/Q VGND VGND VPWR VPWR _20148_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22727__B1 _21121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11944__A _11934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _12783_/Y _12969_/X _12875_/X VGND VGND VPWR VPWR _12970_/Y sky130_fd_sc_hd__a21oi_4
X_20079_ _20079_/A _20079_/B _20079_/C _20079_/D VGND VGND VPWR VPWR _20079_/X sky130_fd_sc_hd__or4_4
X_24956_ _24337_/CLK _15490_/X HRESETn VGND VGND VPWR VPWR _24956_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21137__B _21351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16406__B1 _16315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11921_ _11887_/B _11910_/X _11920_/Y VGND VGND VPWR VPWR _11921_/Y sky130_fd_sc_hd__o21ai_4
X_23907_ _24214_/CLK _23907_/D VGND VGND VPWR VPWR _23907_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24887_ _24889_/CLK _15731_/X HRESETn VGND VGND VPWR VPWR _12536_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14640_ _14632_/X _14639_/Y _25086_/Q _14631_/Y VGND VGND VPWR VPWR _14640_/X sky130_fd_sc_hd__a2bb2o_4
X_11852_ _11849_/Y _11845_/X _11851_/X _11845_/X VGND VGND VPWR VPWR _25530_/D sky130_fd_sc_hd__a2bb2o_4
X_23838_ _24101_/CLK _19185_/X VGND VGND VPWR VPWR _19183_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _13582_/Y _14571_/B VGND VGND VPWR VPWR _14613_/B sky130_fd_sc_hd__or2_4
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ HWDATA[22] VGND VGND VPWR VPWR _11783_/X sky130_fd_sc_hd__buf_2
X_23769_ _23768_/CLK _23769_/D VGND VGND VPWR VPWR _19376_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__13640__B1 _13639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ _16308_/Y _16305_/X _16309_/X _16305_/X VGND VGND VPWR VPWR _24642_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ _13520_/Y _13516_/X _11867_/X _13521_/X VGND VGND VPWR VPWR _13522_/X sky130_fd_sc_hd__a2bb2o_4
X_25508_ _23717_/CLK _25508_/D HRESETn VGND VGND VPWR VPWR _19900_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17290_ _17289_/X VGND VGND VPWR VPWR _24374_/D sky130_fd_sc_hd__inv_2
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16241_ _16241_/A VGND VGND VPWR VPWR _16241_/X sky130_fd_sc_hd__buf_2
X_13453_ _13421_/A _13453_/B VGND VGND VPWR VPWR _13454_/C sky130_fd_sc_hd__or2_4
X_25439_ _25454_/CLK _25439_/D HRESETn VGND VGND VPWR VPWR _25439_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15932__A2 _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12404_ _12275_/Y _12401_/X _12395_/Y _12403_/X VGND VGND VPWR VPWR _12405_/A sky130_fd_sc_hd__a211o_4
X_16172_ _16171_/Y _16167_/X _15995_/X _16167_/X VGND VGND VPWR VPWR _24688_/D sky130_fd_sc_hd__a2bb2o_4
X_13384_ _13416_/A _13384_/B _13383_/X VGND VGND VPWR VPWR _13384_/X sky130_fd_sc_hd__or3_4
XANTENNA__21600__B _22575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15123_ _24983_/Q VGND VGND VPWR VPWR _15424_/A sky130_fd_sc_hd__inv_2
XFILLER_126_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12335_ _12335_/A _12335_/B _12335_/C _12334_/X VGND VGND VPWR VPWR _12349_/C sky130_fd_sc_hd__or4_4
XFILLER_154_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15054_ _15053_/X _22713_/A _15053_/X _22713_/A VGND VGND VPWR VPWR _15054_/X sky130_fd_sc_hd__a2bb2o_4
X_19931_ _19925_/Y VGND VGND VPWR VPWR _19931_/X sky130_fd_sc_hd__buf_2
X_12266_ _24773_/Q VGND VGND VPWR VPWR _12266_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22712__A _16427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ _13999_/C VGND VGND VPWR VPWR _14015_/B sky130_fd_sc_hd__inv_2
X_19862_ _19861_/Y VGND VGND VPWR VPWR _19862_/X sky130_fd_sc_hd__buf_2
XANTENNA__20201__A2_N _20198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17806__A _17752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12197_ _12197_/A VGND VGND VPWR VPWR _12197_/X sky130_fd_sc_hd__buf_2
X_18813_ _18810_/A _18810_/B VGND VGND VPWR VPWR _18813_/Y sky130_fd_sc_hd__nand2_4
X_19793_ _16870_/X VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__buf_2
XFILLER_110_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22718__B1 _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11854__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18744_ _18744_/A _18744_/B VGND VGND VPWR VPWR _18745_/C sky130_fd_sc_hd__or2_4
XFILLER_83_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15956_ _15938_/X _15943_/X HWDATA[25] _24778_/Q _15941_/X VGND VGND VPWR VPWR _24778_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12131__B1 _11871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14907_ _14906_/Y VGND VGND VPWR VPWR _15231_/A sky130_fd_sc_hd__buf_2
X_15887_ _15880_/A VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__buf_2
X_18675_ _18643_/X _18674_/X VGND VGND VPWR VPWR _18713_/A sky130_fd_sc_hd__or2_4
XFILLER_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18637__A _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17626_ _17520_/Y _17626_/B VGND VGND VPWR VPWR _17626_/Y sky130_fd_sc_hd__nand2_4
X_14838_ _14840_/A _14836_/X _14235_/Y _14837_/X VGND VGND VPWR VPWR _14838_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14769_ _14769_/A VGND VGND VPWR VPWR _14769_/X sky130_fd_sc_hd__buf_2
X_17557_ _11754_/Y _24326_/Q _11754_/Y _24326_/Q VGND VGND VPWR VPWR _17560_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19898__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16157__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _16533_/A VGND VGND VPWR VPWR _16508_/X sky130_fd_sc_hd__buf_2
X_17488_ _17487_/Y VGND VGND VPWR VPWR _18361_/A sky130_fd_sc_hd__buf_2
XANTENNA__24903__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19227_ _19224_/Y _19225_/X _19226_/X _19225_/X VGND VGND VPWR VPWR _23823_/D sky130_fd_sc_hd__a2bb2o_4
X_16439_ _15121_/Y _16435_/X _16153_/X _16438_/X VGND VGND VPWR VPWR _16439_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_212_0_HCLK clkbuf_7_106_0_HCLK/X VGND VGND VPWR VPWR _24430_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_164_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19158_ _19158_/A VGND VGND VPWR VPWR _19158_/Y sky130_fd_sc_hd__inv_2
X_18109_ _17973_/X _18108_/X _24251_/Q _18031_/X VGND VGND VPWR VPWR _24251_/D sky130_fd_sc_hd__o22a_4
XFILLER_173_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19089_ _23871_/Q VGND VGND VPWR VPWR _19089_/Y sky130_fd_sc_hd__inv_2
X_21120_ _21040_/Y VGND VGND VPWR VPWR _21121_/A sky130_fd_sc_hd__buf_2
XANTENNA__11748__B _22694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21051_ _12613_/A _15662_/Y _21049_/X _21050_/X VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__a211o_4
XFILLER_207_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18625__A1 _24538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22979__D _22978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16620__A _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20002_ _20002_/A VGND VGND VPWR VPWR _21822_/B sky130_fd_sc_hd__inv_2
XANTENNA__21238__A _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23156__C _23151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24810_ _24812_/CLK _24810_/D HRESETn VGND VGND VPWR VPWR _24810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_228_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19931__A _19925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15163__A2_N _24588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24741_ _24372_/CLK _24741_/D HRESETn VGND VGND VPWR VPWR _24741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21953_ _21476_/A _21953_/B VGND VGND VPWR VPWR _21953_/X sky130_fd_sc_hd__or2_4
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20904_ _20904_/A VGND VGND VPWR VPWR _20904_/X sky130_fd_sc_hd__buf_2
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17451__A _13818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24672_ _24552_/CLK _16225_/X HRESETn VGND VGND VPWR VPWR _16224_/A sky130_fd_sc_hd__dfrtp_4
X_21884_ _11728_/X VGND VGND VPWR VPWR _22443_/A sky130_fd_sc_hd__buf_2
XFILLER_243_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23134__B1 _12899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _24295_/CLK _23623_/D VGND VGND VPWR VPWR _19805_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20842_/A VGND VGND VPWR VPWR _20836_/A sky130_fd_sc_hd__buf_2
XFILLER_70_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22342__D1 _22341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23554_ _23553_/CLK _23554_/D VGND VGND VPWR VPWR _23554_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20766_ _20761_/X _20764_/Y _15608_/A _20765_/X VGND VGND VPWR VPWR _20766_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24644__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _22493_/X _22500_/Y _22501_/X _22504_/X VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _23400_/CLK _20189_/X VGND VGND VPWR VPWR _20188_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _20724_/A VGND VGND VPWR VPWR _20788_/A sky130_fd_sc_hd__buf_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25224_ _25223_/CLK _14158_/X HRESETn VGND VGND VPWR VPWR _14125_/A sky130_fd_sc_hd__dfrtp_4
X_22436_ _21101_/X VGND VGND VPWR VPWR _22436_/X sky130_fd_sc_hd__buf_2
XFILLER_164_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11936__B1 RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25155_ _24012_/CLK _14401_/X HRESETn VGND VGND VPWR VPWR _20475_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_109_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22367_ _21947_/A _19902_/Y _21209_/A VGND VGND VPWR VPWR _22367_/X sky130_fd_sc_hd__o21a_4
X_12120_ _25479_/Q VGND VGND VPWR VPWR _12120_/Y sky130_fd_sc_hd__inv_2
X_24106_ _23647_/CLK _24106_/D HRESETn VGND VGND VPWR VPWR _24106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21318_ _21307_/B _21312_/X _21314_/X _24722_/Q _21317_/X VGND VGND VPWR VPWR _21318_/X
+ sky130_fd_sc_hd__a32o_4
X_25086_ _23703_/CLK _14640_/X HRESETn VGND VGND VPWR VPWR _25086_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22298_ _22298_/A VGND VGND VPWR VPWR _22298_/X sky130_fd_sc_hd__buf_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22948__B1 _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12051_ _12049_/Y _12050_/X _25494_/Q _12050_/X VGND VGND VPWR VPWR _25495_/D sky130_fd_sc_hd__a2bb2o_4
X_24037_ _24042_/CLK _24037_/D HRESETn VGND VGND VPWR VPWR _13129_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21249_ _21271_/A _20230_/Y VGND VGND VPWR VPWR _21250_/C sky130_fd_sc_hd__or2_4
XFILLER_78_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16530__A _14420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ _12373_/Y _15808_/X _11763_/X _15808_/X VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__a2bb2o_4
X_16790_ HWDATA[4] VGND VGND VPWR VPWR _19085_/A sky130_fd_sc_hd__buf_2
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15850__A1 _15833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15741_ _15726_/X VGND VGND VPWR VPWR _15741_/X sky130_fd_sc_hd__buf_2
XANTENNA__15850__B2 _15802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ _12855_/A _12777_/X _12855_/C _12952_/X VGND VGND VPWR VPWR _12956_/B sky130_fd_sc_hd__or4_4
X_24939_ _23717_/CLK _24939_/D HRESETn VGND VGND VPWR VPWR _11736_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_104_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11904_ _25523_/Q _11902_/Y _11898_/B _11903_/X VGND VGND VPWR VPWR _25523_/D sky130_fd_sc_hd__o22a_4
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14200__D _13786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15672_ _21170_/A VGND VGND VPWR VPWR _15673_/A sky130_fd_sc_hd__inv_2
X_18460_ _18710_/A VGND VGND VPWR VPWR _18493_/A sky130_fd_sc_hd__buf_2
XFILLER_206_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12884_ _12878_/A _12872_/X _12883_/X _12880_/B VGND VGND VPWR VPWR _12885_/A sky130_fd_sc_hd__a211o_4
XPHY_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14622_/Y _13647_/X _25086_/Q _13645_/X VGND VGND VPWR VPWR _14639_/A sky130_fd_sc_hd__o22a_4
X_17411_ _24000_/Q _17409_/A VGND VGND VPWR VPWR _17411_/X sky130_fd_sc_hd__or2_4
XPHY_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11803_/X VGND VGND VPWR VPWR _11835_/X sky130_fd_sc_hd__buf_2
X_18391_ _18379_/A VGND VGND VPWR VPWR _18391_/X sky130_fd_sc_hd__buf_2
XANTENNA__16600__A1_N _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17315_/X _17342_/B _17342_/C VGND VGND VPWR VPWR _24361_/D sky130_fd_sc_hd__and3_4
XFILLER_199_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14058_/X _14554_/C _14063_/Y VGND VGND VPWR VPWR _14555_/B sky130_fd_sc_hd__or4_4
XFILLER_186_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ HWDATA[27] VGND VGND VPWR VPWR _11766_/X sky130_fd_sc_hd__buf_2
XANTENNA__18611__A2_N _18737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _12109_/A _12107_/X _12109_/C _13504_/X VGND VGND VPWR VPWR _13506_/A sky130_fd_sc_hd__or4_4
X_17273_ _24377_/Q VGND VGND VPWR VPWR _17274_/A sky130_fd_sc_hd__inv_2
XFILLER_201_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _14485_/A VGND VGND VPWR VPWR _14485_/X sky130_fd_sc_hd__buf_2
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11687_/X _11697_/B _11693_/X _11697_/D VGND VGND VPWR VPWR _11709_/C sky130_fd_sc_hd__or4_4
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _16224_/A VGND VGND VPWR VPWR _16224_/Y sky130_fd_sc_hd__inv_2
X_19012_ _19151_/A VGND VGND VPWR VPWR _19012_/X sky130_fd_sc_hd__buf_2
X_13436_ _13468_/A _23614_/Q VGND VGND VPWR VPWR _13437_/C sky130_fd_sc_hd__or2_4
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16155_ _16152_/Y _16148_/X _16153_/X _16154_/X VGND VGND VPWR VPWR _24695_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22145__C _22145_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11849__A _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13367_ _13241_/X _13363_/X _13366_/X VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__or3_4
XANTENNA__14225__A _20686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15106_ _25000_/Q _24604_/Q _15305_/A _15105_/Y VGND VGND VPWR VPWR _15116_/A sky130_fd_sc_hd__o22a_4
XFILLER_154_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12318_ _24852_/Q VGND VGND VPWR VPWR _12318_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_42_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _24684_/CLK sky130_fd_sc_hd__clkbuf_1
X_16086_ _11729_/X _15659_/B VGND VGND VPWR VPWR _16086_/X sky130_fd_sc_hd__or2_4
X_13298_ _13254_/X _13295_/X _13297_/X VGND VGND VPWR VPWR _13298_/X sky130_fd_sc_hd__and3_4
XFILLER_108_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15037_ _15037_/A VGND VGND VPWR VPWR _15037_/Y sky130_fd_sc_hd__inv_2
X_19914_ _23584_/Q VGND VGND VPWR VPWR _19914_/Y sky130_fd_sc_hd__inv_2
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12249_ _12239_/X _12242_/X _12245_/X _12249_/D VGND VGND VPWR VPWR _12249_/X sky130_fd_sc_hd__or4_4
XANTENNA__23257__B _23254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21058__A _21058_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _19843_/Y _19839_/X _19796_/X _19844_/X VGND VGND VPWR VPWR _23610_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19776_ _19775_/Y _19773_/X _19728_/X _19773_/X VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16988_ _16065_/A _24385_/Q _16065_/Y _16987_/Y VGND VGND VPWR VPWR _16988_/X sky130_fd_sc_hd__o22a_4
X_18727_ _18703_/A _18727_/B VGND VGND VPWR VPWR _18728_/C sky130_fd_sc_hd__or2_4
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15939_ _15793_/X _15870_/B VGND VGND VPWR VPWR _15939_/X sky130_fd_sc_hd__or2_4
X_18658_ _16594_/Y _18657_/X _16594_/Y _18657_/X VGND VGND VPWR VPWR _18659_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23116__B1 _24850_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17609_ _17663_/A _17609_/B VGND VGND VPWR VPWR _17610_/D sky130_fd_sc_hd__and2_4
XFILLER_212_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18589_ _18568_/X _18588_/X _18598_/C VGND VGND VPWR VPWR _24168_/D sky130_fd_sc_hd__and3_4
X_20620_ _20620_/A VGND VGND VPWR VPWR _20621_/B sky130_fd_sc_hd__buf_2
XANTENNA__21678__B1 _18306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15824__A1_N _12350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21142__A2 _21375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20551_ _20550_/Y VGND VGND VPWR VPWR _20551_/X sky130_fd_sc_hd__buf_2
XFILLER_20_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16615__A _16615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23270_ _20960_/Y _21606_/A _20821_/Y _22298_/A VGND VGND VPWR VPWR _23270_/X sky130_fd_sc_hd__o22a_4
X_20482_ _23978_/Q VGND VGND VPWR VPWR _20503_/B sky130_fd_sc_hd__inv_2
XFILLER_138_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22221_ _22221_/A _22221_/B _22220_/X VGND VGND VPWR VPWR _22221_/X sky130_fd_sc_hd__or3_4
XANTENNA__11759__A _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15839__A1_N _12327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19926__A _19925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18830__A pwm_S7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22152_ _24351_/Q _23093_/A _22810_/A VGND VGND VPWR VPWR _22152_/X sky130_fd_sc_hd__a21o_4
XFILLER_160_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21103_ _21103_/A VGND VGND VPWR VPWR _21104_/B sky130_fd_sc_hd__buf_2
X_22083_ _22390_/A _22080_/X _22083_/C VGND VGND VPWR VPWR _22083_/X sky130_fd_sc_hd__and3_4
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21034_ _21605_/A VGND VGND VPWR VPWR _21034_/X sky130_fd_sc_hd__buf_2
XFILLER_160_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22158__A1 _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22985_ _22985_/A _22985_/B VGND VGND VPWR VPWR _22985_/X sky130_fd_sc_hd__or2_4
XFILLER_28_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13843__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20600__A _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24896__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24724_ _24726_/CLK _16079_/X HRESETn VGND VGND VPWR VPWR _16078_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_227_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21936_ _21936_/A VGND VGND VPWR VPWR _21941_/A sky130_fd_sc_hd__buf_2
XFILLER_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24825__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24655_ _24194_/CLK _24655_/D HRESETn VGND VGND VPWR VPWR _24655_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21867_ _21731_/A _21863_/X _21866_/X VGND VGND VPWR VPWR _21867_/Y sky130_fd_sc_hd__o21ai_4
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23597_/CLK _19854_/X VGND VGND VPWR VPWR _19853_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _20818_/A _20818_/B VGND VGND VPWR VPWR _20818_/X sky130_fd_sc_hd__and2_4
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24586_ _24592_/CLK _24586_/D HRESETn VGND VGND VPWR VPWR _15134_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21798_ _22549_/B _21797_/X _13581_/Y _22549_/B VGND VGND VPWR VPWR _21798_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _23560_/CLK _23537_/D VGND VGND VPWR VPWR _23537_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ _13141_/X VGND VGND VPWR VPWR _20749_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14270_/A VGND VGND VPWR VPWR _14270_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23468_ _23794_/CLK _23468_/D VGND VGND VPWR VPWR _20232_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_7_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _13271_/A VGND VGND VPWR VPWR _13320_/A sky130_fd_sc_hd__buf_2
X_25207_ _25204_/CLK _14226_/X HRESETn VGND VGND VPWR VPWR _20686_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22419_ _22283_/X _22418_/X _22148_/C _24832_/Q _22286_/X VGND VGND VPWR VPWR _22419_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22633__A2 _21320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23399_ _23400_/CLK _23399_/D VGND VGND VPWR VPWR _23399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16848__B1 _11830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13152_ _13306_/A VGND VGND VPWR VPWR _13285_/A sky130_fd_sc_hd__buf_2
X_25138_ _25215_/CLK _25138_/D HRESETn VGND VGND VPWR VPWR _14455_/A sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_1_0_HCLK clkbuf_7_0_0_HCLK/X VGND VGND VPWR VPWR _23408_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_29_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_58_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12103_ _12102_/X VGND VGND VPWR VPWR _12109_/A sky130_fd_sc_hd__buf_2
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13083_ _13083_/A _13083_/B VGND VGND VPWR VPWR _13085_/B sky130_fd_sc_hd__or2_4
X_17960_ _17945_/A _17958_/X _17960_/C VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__and3_4
X_25069_ _25066_/CLK _14756_/X HRESETn VGND VGND VPWR VPWR _14723_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12034_ _12032_/Y _20977_/A _12032_/Y _20977_/A VGND VGND VPWR VPWR _12034_/X sky130_fd_sc_hd__a2bb2o_4
X_16911_ _22994_/A _17824_/A _23205_/A _16910_/Y VGND VGND VPWR VPWR _16911_/X sky130_fd_sc_hd__a2bb2o_4
X_17891_ _16929_/Y _17891_/B VGND VGND VPWR VPWR _17892_/C sky130_fd_sc_hd__nand2_4
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23175__A1_N _17245_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19630_ _19628_/Y _19625_/X _19629_/X _19625_/X VGND VGND VPWR VPWR _23683_/D sky130_fd_sc_hd__a2bb2o_4
X_16842_ _16841_/Y _16839_/X _15756_/X _16839_/X VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22149__A1 _21714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19561_ _19559_/Y _19557_/X _19560_/X _19557_/X VGND VGND VPWR VPWR _23705_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21606__A _21606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13985_ _23941_/Q VGND VGND VPWR VPWR _13985_/X sky130_fd_sc_hd__buf_2
X_16773_ _16782_/A VGND VGND VPWR VPWR _16773_/X sky130_fd_sc_hd__buf_2
XANTENNA__18187__A _18059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18512_ _18486_/X _18503_/X _18487_/A VGND VGND VPWR VPWR _18512_/X sky130_fd_sc_hd__o21a_4
XFILLER_207_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12936_ _12912_/A _12933_/X VGND VGND VPWR VPWR _12936_/X sky130_fd_sc_hd__or2_4
X_15724_ _15557_/X _15722_/X _15723_/X _24890_/Q _15720_/X VGND VGND VPWR VPWR _15724_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_74_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19492_ _21959_/B _19489_/X _11952_/X _19489_/X VGND VGND VPWR VPWR _19492_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24566__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18443_ _18443_/A _18443_/B _18443_/C _18443_/D VGND VGND VPWR VPWR _18457_/B sky130_fd_sc_hd__or4_4
XFILLER_179_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12867_ _12869_/B VGND VGND VPWR VPWR _12868_/B sky130_fd_sc_hd__inv_2
X_15655_ _21299_/A VGND VGND VPWR VPWR _15655_/X sky130_fd_sc_hd__buf_2
XFILLER_221_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15587__B1 _11776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _16245_/A VGND VGND VPWR VPWR _11818_/X sky130_fd_sc_hd__buf_2
X_14606_ _14575_/X _14595_/X _14605_/Y _14599_/X _14568_/A VGND VGND VPWR VPWR _25095_/D
+ sky130_fd_sc_hd__a32o_4
X_15586_ _15586_/A VGND VGND VPWR VPWR _15586_/Y sky130_fd_sc_hd__inv_2
X_18374_ _18372_/A VGND VGND VPWR VPWR _18374_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22857__C1 _22856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17328__A1 _17263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12798_ _25375_/Q _21537_/A _12796_/Y _12797_/Y VGND VGND VPWR VPWR _12798_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22321__B2 _21375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _21560_/A _14519_/X _21352_/A _14514_/X VGND VGND VPWR VPWR _14537_/X sky130_fd_sc_hd__o22a_4
X_17325_ _17324_/X VGND VGND VPWR VPWR _24366_/D sky130_fd_sc_hd__inv_2
X_11749_ _11749_/A VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__buf_2
XFILLER_175_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12963__A _12793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ _14468_/A VGND VGND VPWR VPWR _14468_/X sky130_fd_sc_hd__buf_2
X_17256_ _17197_/Y _17178_/A _17252_/X _17256_/D VGND VGND VPWR VPWR _17256_/X sky130_fd_sc_hd__or4_4
XFILLER_174_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13419_ _13451_/A _13417_/X _13419_/C VGND VGND VPWR VPWR _13423_/B sky130_fd_sc_hd__and3_4
X_16207_ _23218_/A VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
X_17187_ _17293_/A VGND VGND VPWR VPWR _17294_/A sky130_fd_sc_hd__inv_2
XFILLER_162_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14399_ _20475_/C VGND VGND VPWR VPWR _20514_/D sky130_fd_sc_hd__inv_2
XFILLER_128_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16138_ _22763_/A VGND VGND VPWR VPWR _16138_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17500__B2 _17499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _16044_/A VGND VGND VPWR VPWR _16069_/X sky130_fd_sc_hd__buf_2
XANTENNA__17266__A _17266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15511__B1 HADDR[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20399__B1 _19643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22900__A _22944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20938__A2 _20854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19828_ _23615_/Q VGND VGND VPWR VPWR _19828_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23337__B1 _22479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19759_ _19758_/Y _19756_/X _19692_/X _19756_/X VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18097__A _18097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22770_ _22769_/X VGND VGND VPWR VPWR _22770_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22560__A1 _16606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21721_ _21542_/X _21717_/Y _22723_/A _21720_/X VGND VGND VPWR VPWR _21721_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15578__B1 _11763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24440_ _24437_/CLK _16826_/X HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
X_21652_ _21632_/X _21651_/X _21511_/X VGND VGND VPWR VPWR _21652_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_178_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20603_ _14103_/A _20603_/B _20603_/C VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__and3_4
X_24371_ _24641_/CLK _24371_/D HRESETn VGND VGND VPWR VPWR _24371_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21583_ _21577_/A _21583_/B VGND VGND VPWR VPWR _21583_/X sky130_fd_sc_hd__or2_4
XFILLER_193_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22863__A2 _22530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23322_ _24821_/Q _23322_/B VGND VGND VPWR VPWR _23322_/X sky130_fd_sc_hd__or2_4
XFILLER_166_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20534_ _20534_/A VGND VGND VPWR VPWR _20534_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22337__A1_N _14816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23253_ _23253_/A _23253_/B _23253_/C VGND VGND VPWR VPWR _23253_/X sky130_fd_sc_hd__and3_4
XANTENNA__19656__A _19148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20465_ _20448_/X _20457_/X VGND VGND VPWR VPWR _20465_/X sky130_fd_sc_hd__and2_4
XANTENNA__15750__B1 _24876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22204_ _22204_/A _22199_/X _22204_/C VGND VGND VPWR VPWR _22204_/X sky130_fd_sc_hd__and3_4
XFILLER_192_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23184_ _22897_/A VGND VGND VPWR VPWR _23184_/X sky130_fd_sc_hd__buf_2
X_20396_ _21818_/B _20391_/X _19639_/A _20391_/X VGND VGND VPWR VPWR _23407_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22135_ _22129_/X _22131_/Y _22133_/Y _22134_/X _21565_/Y VGND VGND VPWR VPWR _22135_/X
+ sky130_fd_sc_hd__o41a_4
XANTENNA__15502__B1 HADDR[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22066_ _22066_/A VGND VGND VPWR VPWR _22066_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23040__A2 _23031_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22810__A _22810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21051__A1 _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21017_ _23980_/Q _23981_/Q _21018_/B VGND VGND VPWR VPWR _23980_/D sky130_fd_sc_hd__o21a_4
XFILLER_248_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21426__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13816__B1 _13524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11952__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ _25284_/Q VGND VGND VPWR VPWR _13770_/X sky130_fd_sc_hd__buf_2
XFILLER_216_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22968_ _24471_/Q _22968_/B _22853_/X VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__and3_4
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22551__A1 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12721_ _12623_/D _12718_/B VGND VGND VPWR VPWR _12722_/C sky130_fd_sc_hd__nand2_4
XFILLER_243_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21919_ _22235_/A _21919_/B _21918_/X VGND VGND VPWR VPWR _21919_/X sky130_fd_sc_hd__and3_4
X_24707_ _25444_/CLK _24707_/D HRESETn VGND VGND VPWR VPWR _22994_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_15_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22899_ _24538_/Q _21085_/A _22815_/X _22898_/X VGND VGND VPWR VPWR _22900_/C sky130_fd_sc_hd__a211o_4
XFILLER_188_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15440_ _15439_/X VGND VGND VPWR VPWR _15440_/X sky130_fd_sc_hd__buf_2
X_12652_ _12654_/B VGND VGND VPWR VPWR _12657_/B sky130_fd_sc_hd__inv_2
X_24638_ _24629_/CLK _16321_/X HRESETn VGND VGND VPWR VPWR _24638_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14241__B1 _13806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18658__A1_N _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21161__A _21161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _15376_/A _15306_/B _15380_/A _15384_/B VGND VGND VPWR VPWR _15377_/B sky130_fd_sc_hd__or4_4
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12583_/A VGND VGND VPWR VPWR _12619_/B sky130_fd_sc_hd__inv_2
X_24569_ _24602_/CLK _16505_/X HRESETn VGND VGND VPWR VPWR _24569_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12783__A _25380_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _25181_/Q _14311_/X _25180_/Q _14316_/X VGND VGND VPWR VPWR _14322_/X sky130_fd_sc_hd__o22a_4
X_17110_ _17042_/C _17110_/B VGND VGND VPWR VPWR _17120_/B sky130_fd_sc_hd__or2_4
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18090_ _18090_/A _18090_/B VGND VGND VPWR VPWR _18092_/B sky130_fd_sc_hd__or2_4
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17041_/A VGND VGND VPWR VPWR _17042_/D sky130_fd_sc_hd__inv_2
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _13958_/A _13924_/B _13924_/C _14252_/Y VGND VGND VPWR VPWR _14254_/B sky130_fd_sc_hd__and4_4
XFILLER_183_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19566__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _11993_/Y _13203_/Y _11985_/A VGND VGND VPWR VPWR _13267_/A sky130_fd_sc_hd__o21a_4
X_14184_ _14178_/Y _14119_/X _14120_/X _14183_/X VGND VGND VPWR VPWR _14185_/A sky130_fd_sc_hd__o22a_4
XFILLER_152_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13135_ _13135_/A _13134_/X VGND VGND VPWR VPWR _13136_/B sky130_fd_sc_hd__or2_4
XANTENNA__17086__A _17074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18992_ _14674_/A VGND VGND VPWR VPWR _18992_/X sky130_fd_sc_hd__buf_2
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13066_ _12312_/X _13066_/B VGND VGND VPWR VPWR _13066_/X sky130_fd_sc_hd__or2_4
X_17943_ _17943_/A _17943_/B VGND VGND VPWR VPWR _17945_/B sky130_fd_sc_hd__or2_4
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_116_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24867_/CLK sky130_fd_sc_hd__clkbuf_1
X_12017_ _12002_/X VGND VGND VPWR VPWR _12017_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17874_ _17861_/B _17861_/D _17798_/X _17871_/B VGND VGND VPWR VPWR _17875_/A sky130_fd_sc_hd__a211o_4
XFILLER_66_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_179_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _24112_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19613_ _19611_/Y _19606_/X _19612_/X _19606_/X VGND VGND VPWR VPWR _23688_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22790__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24747__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16825_ _16810_/X VGND VGND VPWR VPWR _16825_/X sky130_fd_sc_hd__buf_2
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13807__B1 _13806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12958__A _12855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11862__A _14412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19544_ _21502_/B _19541_/X _11964_/X _19541_/X VGND VGND VPWR VPWR _23710_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16756_ _23037_/A VGND VGND VPWR VPWR _16756_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13968_ _13967_/X VGND VGND VPWR VPWR _13968_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14480__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21345__A2 _22610_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15707_ _14629_/B _15703_/X VGND VGND VPWR VPWR _15707_/X sky130_fd_sc_hd__and2_4
XFILLER_206_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12919_ _12834_/Y _12913_/X _12883_/X _12915_/Y VGND VGND VPWR VPWR _12920_/A sky130_fd_sc_hd__a211o_4
X_19475_ _18184_/B VGND VGND VPWR VPWR _19475_/Y sky130_fd_sc_hd__inv_2
X_13899_ _24979_/Q _24978_/Q _13899_/C VGND VGND VPWR VPWR _13899_/X sky130_fd_sc_hd__or3_4
X_16687_ _24501_/Q VGND VGND VPWR VPWR _16687_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12192__A1_N _25444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18426_ _16273_/A _24165_/Q _16273_/Y _18425_/Y VGND VGND VPWR VPWR _18429_/C sky130_fd_sc_hd__o22a_4
XFILLER_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15638_ _24902_/Q VGND VGND VPWR VPWR _15638_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22167__A _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18357_ _18357_/A VGND VGND VPWR VPWR _18357_/Y sky130_fd_sc_hd__inv_2
X_15569_ _15569_/A VGND VGND VPWR VPWR _15589_/A sky130_fd_sc_hd__inv_2
XFILLER_203_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17308_ _17308_/A VGND VGND VPWR VPWR _24370_/D sky130_fd_sc_hd__inv_2
XFILLER_148_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18288_ _17712_/A VGND VGND VPWR VPWR _18288_/X sky130_fd_sc_hd__buf_2
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23067__A1_N _17266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17239_ _17239_/A _17239_/B _17233_/X _17239_/D VGND VGND VPWR VPWR _17240_/B sky130_fd_sc_hd__or4_4
XFILLER_163_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20250_ _20247_/Y _20248_/X _20249_/X _20248_/X VGND VGND VPWR VPWR _20250_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23270__A2 _21606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20181_ _23488_/Q VGND VGND VPWR VPWR _20181_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_75_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23940_ _25106_/CLK _23940_/D HRESETn VGND VGND VPWR VPWR _23940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_215_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23871_ _23871_/CLK _19092_/X VGND VGND VPWR VPWR _23871_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12868__A _25404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22822_ _24536_/Q _22541_/A _22542_/A _22821_/X VGND VGND VPWR VPWR _22822_/X sky130_fd_sc_hd__a211o_4
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14471__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21336__A2 _21312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25541_ _25539_/CLK _25541_/D HRESETn VGND VGND VPWR VPWR _11802_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22753_ _16594_/A _21067_/X _21755_/A _22752_/X VGND VGND VPWR VPWR _22754_/C sky130_fd_sc_hd__a211o_4
XFILLER_198_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21887__A3 _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24070__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21704_ _21704_/A _21660_/X VGND VGND VPWR VPWR _21704_/Y sky130_fd_sc_hd__nor2_4
XFILLER_213_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25472_ _25215_/CLK _12179_/X HRESETn VGND VGND VPWR VPWR SCLK_S3 sky130_fd_sc_hd__dfstp_4
X_22684_ _16515_/Y _22684_/B VGND VGND VPWR VPWR _22684_/X sky130_fd_sc_hd__and2_4
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24423_ _24425_/CLK _24423_/D HRESETn VGND VGND VPWR VPWR _24423_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21635_ _21259_/A VGND VGND VPWR VPWR _22090_/A sky130_fd_sc_hd__buf_2
XFILLER_139_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15971__B1 _15970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16075__A _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19162__B1 _19048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24354_ _24354_/CLK _17373_/Y HRESETn VGND VGND VPWR VPWR _17193_/A sky130_fd_sc_hd__dfrtp_4
X_21566_ _14279_/Y _21375_/X VGND VGND VPWR VPWR _21566_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23305_ _23137_/X _23303_/X _23139_/X _23304_/X VGND VGND VPWR VPWR _23306_/B sky130_fd_sc_hd__o22a_4
XFILLER_165_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20517_ _24014_/Q _20456_/X _20478_/B VGND VGND VPWR VPWR _24014_/D sky130_fd_sc_hd__a21o_4
X_24285_ _24272_/CLK _17816_/Y HRESETn VGND VGND VPWR VPWR _24285_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21497_ _21497_/A _21497_/B VGND VGND VPWR VPWR _21497_/X sky130_fd_sc_hd__or2_4
XANTENNA__12108__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23236_ _23236_/A VGND VGND VPWR VPWR _23236_/Y sky130_fd_sc_hd__inv_2
X_20448_ _24098_/Q VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__buf_2
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11947__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23167_ _23167_/A VGND VGND VPWR VPWR _23167_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20379_ _20379_/A VGND VGND VPWR VPWR _21480_/B sky130_fd_sc_hd__inv_2
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22118_ _14489_/Y _21375_/X _25112_/Q _22129_/B VGND VGND VPWR VPWR _22118_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23098_ _21427_/A _23096_/Y _22844_/X _23097_/X VGND VGND VPWR VPWR _23099_/A sky130_fd_sc_hd__o22a_4
XANTENNA__20979__B _12168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17228__B1 _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14940_ _15188_/A _14939_/A _15182_/A _14939_/Y VGND VGND VPWR VPWR _14940_/X sky130_fd_sc_hd__o22a_4
X_22049_ _22036_/A _22045_/X _22046_/X _22047_/X _22048_/X VGND VGND VPWR VPWR _22049_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17634__A _17691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18976__B1 _18975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24840__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14871_ _14837_/X _14870_/X _15479_/A _14840_/A VGND VGND VPWR VPWR _14871_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16618_/A VGND VGND VPWR VPWR _16610_/X sky130_fd_sc_hd__buf_2
XFILLER_217_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13822_ _13822_/A _13822_/B VGND VGND VPWR VPWR _14462_/A sky130_fd_sc_hd__or2_4
X_17590_ _17667_/A _17581_/Y _17589_/X VGND VGND VPWR VPWR _17590_/X sky130_fd_sc_hd__or3_4
XFILLER_232_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13753_ _14769_/A _13748_/X _14789_/A _13597_/X VGND VGND VPWR VPWR _13753_/X sky130_fd_sc_hd__or4_4
X_16541_ _16539_/Y _16533_/X _16364_/X _16540_/X VGND VGND VPWR VPWR _24556_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12704_ _12704_/A VGND VGND VPWR VPWR _12705_/B sky130_fd_sc_hd__inv_2
X_19260_ _22372_/B _19259_/X _16872_/X _19259_/X VGND VGND VPWR VPWR _19260_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23090__B _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13684_ _13652_/A _25302_/Q _25303_/Q VGND VGND VPWR VPWR _13684_/X sky130_fd_sc_hd__a21o_4
X_16472_ _16472_/A VGND VGND VPWR VPWR _16472_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18211_ _17991_/X _18211_/B _18211_/C VGND VGND VPWR VPWR _18212_/C sky130_fd_sc_hd__and3_4
XFILLER_231_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12635_ _12521_/Y _12633_/A VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__or2_4
X_15423_ _15423_/A _15423_/B VGND VGND VPWR VPWR _15424_/B sky130_fd_sc_hd__or2_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19191_ _19196_/A VGND VGND VPWR VPWR _19191_/X sky130_fd_sc_hd__buf_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13402__A _13217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15354_ _15354_/A _15357_/B VGND VGND VPWR VPWR _15355_/C sky130_fd_sc_hd__or2_4
X_18142_ _18072_/X _18142_/B VGND VGND VPWR VPWR _18142_/X sky130_fd_sc_hd__or2_4
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12566_ _12566_/A _12566_/B _12566_/C _12565_/X VGND VGND VPWR VPWR _12566_/X sky130_fd_sc_hd__or4_4
XFILLER_200_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22715__A _21879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ _14305_/A _14316_/A VGND VGND VPWR VPWR _14305_/X sky130_fd_sc_hd__or2_4
XFILLER_172_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _15285_/A VGND VGND VPWR VPWR _25017_/D sky130_fd_sc_hd__inv_2
X_18073_ _18072_/X _19376_/A VGND VGND VPWR VPWR _18073_/X sky130_fd_sc_hd__or2_4
X_12497_ _12278_/Y _12500_/B VGND VGND VPWR VPWR _12501_/B sky130_fd_sc_hd__or2_4
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14236_ _14235_/Y _14233_/X _13846_/X _14233_/X VGND VGND VPWR VPWR _25205_/D sky130_fd_sc_hd__a2bb2o_4
X_17024_ _16068_/Y _24384_/Q _16078_/Y _24381_/Q VGND VGND VPWR VPWR _17024_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14234__A1_N _14227_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23252__A2 _22485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11857__A _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ _14153_/X _14166_/Y _25221_/Q _14153_/X VGND VGND VPWR VPWR _14167_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13118_ _12387_/X _13121_/A VGND VGND VPWR VPWR _13118_/X sky130_fd_sc_hd__or2_4
XANTENNA__24928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14098_ _14082_/A VGND VGND VPWR VPWR _20549_/B sky130_fd_sc_hd__buf_2
X_18975_ _19091_/A VGND VGND VPWR VPWR _18975_/X sky130_fd_sc_hd__buf_2
X_13049_ _13049_/A _13046_/B _13049_/C VGND VGND VPWR VPWR _13049_/X sky130_fd_sc_hd__or3_4
X_17926_ _17925_/Y _15922_/A _17924_/B VGND VGND VPWR VPWR _17926_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23265__B _22954_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18967__B1 _17433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24581__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21066__A _21066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _17757_/D _17562_/X VGND VGND VPWR VPWR _17858_/B sky130_fd_sc_hd__or2_4
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16808_ _24449_/Q VGND VGND VPWR VPWR _16808_/Y sky130_fd_sc_hd__inv_2
X_17788_ _16925_/Y _17788_/B VGND VGND VPWR VPWR _17789_/C sky130_fd_sc_hd__or2_4
XANTENNA__21318__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19527_ _18283_/X _18294_/X _19527_/C _20015_/B VGND VGND VPWR VPWR _19527_/X sky130_fd_sc_hd__or4_4
X_16739_ _16738_/X VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__buf_2
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ _17965_/B VGND VGND VPWR VPWR _19458_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18409_ _24673_/Q _18534_/A _23218_/A _18510_/A VGND VGND VPWR VPWR _18411_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19389_ _17956_/B VGND VGND VPWR VPWR _19389_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22818__A2 _21085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21420_ _21416_/X _21419_/X _14692_/A VGND VGND VPWR VPWR _21420_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12231__A2 _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22625__A _22592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19695__B2 _19675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21351_ _21351_/A VGND VGND VPWR VPWR _22190_/B sky130_fd_sc_hd__buf_2
XANTENNA__15705__B1 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20302_ _20302_/A VGND VGND VPWR VPWR _20302_/Y sky130_fd_sc_hd__inv_2
X_24070_ _24503_/CLK _20939_/Y HRESETn VGND VGND VPWR VPWR _24070_/Q sky130_fd_sc_hd__dfrtp_4
X_21282_ _18268_/A VGND VGND VPWR VPWR _21282_/X sky130_fd_sc_hd__buf_2
X_23021_ _22997_/X _23001_/X _23005_/Y _23020_/X VGND VGND VPWR VPWR HRDATA[21] sky130_fd_sc_hd__a211o_4
X_20233_ _13626_/A _19436_/B _14665_/Y _19346_/B VGND VGND VPWR VPWR _20233_/X sky130_fd_sc_hd__or4_4
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24669__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20164_ _21647_/B _20163_/X _20119_/X _20163_/X VGND VGND VPWR VPWR _23495_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22203__B1 _21121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20095_ _20095_/A VGND VGND VPWR VPWR _20095_/Y sky130_fd_sc_hd__inv_2
X_24972_ _24975_/CLK _24972_/D HRESETn VGND VGND VPWR VPWR _13952_/C sky130_fd_sc_hd__dfrtp_4
X_23923_ _25491_/CLK _23923_/D VGND VGND VPWR VPWR _18942_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_162_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23850_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_242_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23854_ _23871_/CLK _19137_/X VGND VGND VPWR VPWR _13411_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_19_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _23534_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15787__A3 _15782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22805_ _22805_/A _22891_/B VGND VGND VPWR VPWR _22805_/X sky130_fd_sc_hd__and2_4
XFILLER_214_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21704__A _21704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23785_ _24252_/CLK _19334_/X VGND VGND VPWR VPWR _23785_/Q sky130_fd_sc_hd__dfxtp_4
X_20997_ _20997_/A VGND VGND VPWR VPWR _23944_/D sky130_fd_sc_hd__inv_2
XFILLER_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22736_ _22294_/A _22735_/X VGND VGND VPWR VPWR _22736_/Y sky130_fd_sc_hd__nor2_4
X_25524_ _25520_/CLK _25524_/D HRESETn VGND VGND VPWR VPWR _25524_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25455_ _25443_/CLK _25455_/D HRESETn VGND VGND VPWR VPWR _12255_/A sky130_fd_sc_hd__dfrtp_4
X_22667_ _21082_/X _22666_/X VGND VGND VPWR VPWR _22676_/C sky130_fd_sc_hd__and2_4
XANTENNA__19135__B1 _19091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12420_ _12299_/B _12400_/B _12299_/A VGND VGND VPWR VPWR _12421_/C sky130_fd_sc_hd__o21a_4
X_24406_ _24406_/CLK _24406_/D HRESETn VGND VGND VPWR VPWR _24406_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13222__A _13320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21618_ _21412_/A VGND VGND VPWR VPWR _22235_/A sky130_fd_sc_hd__buf_2
X_25386_ _25392_/CLK _25386_/D HRESETn VGND VGND VPWR VPWR _25386_/Q sky130_fd_sc_hd__dfrtp_4
X_22598_ _17362_/A _22677_/B _22597_/X VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__o21a_4
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12351_ _12351_/A VGND VGND VPWR VPWR _12351_/Y sky130_fd_sc_hd__inv_2
X_24337_ _24337_/CLK _17431_/X HRESETn VGND VGND VPWR VPWR _17429_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_194_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21549_ _24619_/Q _21719_/B VGND VGND VPWR VPWR _21549_/X sky130_fd_sc_hd__or2_4
XFILLER_5_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15070_ _15070_/A _15275_/A _15258_/A _14916_/Y VGND VGND VPWR VPWR _15073_/C sky130_fd_sc_hd__or4_4
XFILLER_5_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12282_ _12282_/A _12281_/X VGND VGND VPWR VPWR _12282_/X sky130_fd_sc_hd__or2_4
X_24268_ _24715_/CLK _24268_/D HRESETn VGND VGND VPWR VPWR _16937_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14021_ _14062_/A _14021_/B _14020_/Y _14021_/D VGND VGND VPWR VPWR _14022_/B sky130_fd_sc_hd__or4_4
X_23219_ _24579_/Q _23184_/X _23148_/X VGND VGND VPWR VPWR _23219_/X sky130_fd_sc_hd__o21a_4
XFILLER_107_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19844__A _19838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24199_ _25145_/CLK _18389_/X HRESETn VGND VGND VPWR VPWR _24199_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16121__B1 _15960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17364__A _17364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ _18765_/A _18764_/A _18763_/A _18751_/X VGND VGND VPWR VPWR _18766_/B sky130_fd_sc_hd__or4_4
X_15972_ HWDATA[17] VGND VGND VPWR VPWR _15972_/X sky130_fd_sc_hd__buf_2
XFILLER_110_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17711_ _17711_/A _17711_/B _21704_/A _17711_/D VGND VGND VPWR VPWR _17712_/A sky130_fd_sc_hd__or4_4
X_14923_ _14920_/A _14922_/A _14921_/X _14922_/Y VGND VGND VPWR VPWR _14933_/A sky130_fd_sc_hd__o22a_4
X_18691_ _18630_/Y _18691_/B _18687_/X _18690_/X VGND VGND VPWR VPWR _18700_/A sky130_fd_sc_hd__or4_4
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17642_ _17579_/B _17636_/X _17611_/X _17638_/Y VGND VGND VPWR VPWR _17642_/X sky130_fd_sc_hd__a211o_4
X_14854_ _14840_/A VGND VGND VPWR VPWR _14854_/X sky130_fd_sc_hd__buf_2
XANTENNA__22798__A1_N _17262_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15778__A3 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13805_ _13805_/A VGND VGND VPWR VPWR _13805_/X sky130_fd_sc_hd__buf_2
X_17573_ _17573_/A _17520_/Y VGND VGND VPWR VPWR _17573_/X sky130_fd_sc_hd__or2_4
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11997_ _11663_/B _11986_/X _11996_/Y VGND VGND VPWR VPWR _25501_/D sky130_fd_sc_hd__o21a_4
X_14785_ _14785_/A _14785_/B VGND VGND VPWR VPWR _14785_/X sky130_fd_sc_hd__and2_4
XFILLER_217_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19312_ _19311_/Y _19309_/X _19220_/X _19309_/X VGND VGND VPWR VPWR _19312_/X sky130_fd_sc_hd__a2bb2o_4
X_16524_ _24561_/Q VGND VGND VPWR VPWR _16524_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13736_ _13736_/A _13691_/X VGND VGND VPWR VPWR _13736_/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19243_ _13312_/B VGND VGND VPWR VPWR _19243_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22148__C _22148_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16455_ _16454_/Y _16384_/A _16375_/X _16384_/A VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15935__B1 _24786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13667_ _13667_/A _13667_/B VGND VGND VPWR VPWR _20865_/B sky130_fd_sc_hd__or2_4
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14228__A _14228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15406_ _15082_/Y _15408_/B _15405_/Y VGND VGND VPWR VPWR _15406_/X sky130_fd_sc_hd__o21a_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12618_ _12618_/A _12618_/B _12618_/C _12618_/D VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__or4_4
X_19174_ _19181_/A VGND VGND VPWR VPWR _19174_/X sky130_fd_sc_hd__buf_2
X_13598_ _13597_/X VGND VGND VPWR VPWR _13599_/B sky130_fd_sc_hd__inv_2
X_16386_ _16377_/Y _16384_/X _16385_/X _16384_/X VGND VGND VPWR VPWR _24616_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18125_ _18090_/A _18125_/B VGND VGND VPWR VPWR _18125_/X sky130_fd_sc_hd__or2_4
X_12549_ _25430_/Q _24884_/Q _12616_/B _12548_/Y VGND VGND VPWR VPWR _12549_/X sky130_fd_sc_hd__o22a_4
X_15337_ _15337_/A _15337_/B VGND VGND VPWR VPWR _15340_/B sky130_fd_sc_hd__or2_4
XFILLER_200_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18056_ _18200_/A _23898_/Q VGND VGND VPWR VPWR _18057_/C sky130_fd_sc_hd__or2_4
XANTENNA__24082__D _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ _15268_/A _15259_/X VGND VGND VPWR VPWR _15271_/B sky130_fd_sc_hd__or2_4
XANTENNA__16360__B1 _16070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15163__B2 _15134_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17007_ _17001_/X _17004_/X _17005_/X _17006_/X VGND VGND VPWR VPWR _17007_/X sky130_fd_sc_hd__or4_4
X_14219_ _20675_/A _14207_/B VGND VGND VPWR VPWR _14219_/X sky130_fd_sc_hd__or2_4
XFILLER_99_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22433__B1 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ _14996_/X _15195_/B _15198_/X VGND VGND VPWR VPWR _15199_/X sky130_fd_sc_hd__or3_4
XFILLER_113_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24762__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16112__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17274__A _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18958_ _18958_/A VGND VGND VPWR VPWR _18958_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17909_ _17909_/A VGND VGND VPWR VPWR _17910_/B sky130_fd_sc_hd__inv_2
X_18889_ _18891_/B VGND VGND VPWR VPWR _18890_/A sky130_fd_sc_hd__inv_2
XFILLER_55_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20920_ _13658_/D _20915_/X _20924_/B VGND VGND VPWR VPWR _20920_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__17612__B1 _17611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_235_0_HCLK clkbuf_8_234_0_HCLK/A VGND VGND VPWR VPWR _25106_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12211__A _25446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16966__A2 _16964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20851_ _24051_/Q _13664_/X _20850_/Y VGND VGND VPWR VPWR _20851_/Y sky130_fd_sc_hd__a21oi_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14977__B2 _14976_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16618__A _16618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19365__B1 _19254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23570_ _23560_/CLK _19952_/X VGND VGND VPWR VPWR _23570_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20782_ _22934_/A _20716_/A _20724_/X _20781_/Y VGND VGND VPWR VPWR _20782_/X sky130_fd_sc_hd__o22a_4
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25550__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22521_ _13822_/B _22519_/X _21605_/X _22520_/X VGND VGND VPWR VPWR _22522_/A sky130_fd_sc_hd__o22a_4
XANTENNA__14756__A1_N _14725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25240_ _25105_/CLK _14089_/X HRESETn VGND VGND VPWR VPWR _13999_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_195_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22452_ _22436_/X _22452_/B _22446_/Y _22451_/Y VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__or4_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21403_ _14765_/X _21403_/B VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__or2_4
X_25171_ _25168_/CLK _14345_/X HRESETn VGND VGND VPWR VPWR _25171_/Q sky130_fd_sc_hd__dfrtp_4
X_22383_ _22390_/A _22383_/B _22383_/C VGND VGND VPWR VPWR _22383_/X sky130_fd_sc_hd__and3_4
XFILLER_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24122_ _25145_/CLK _24122_/D HRESETn VGND VGND VPWR VPWR _21002_/A sky130_fd_sc_hd__dfrtp_4
X_21334_ _21591_/A VGND VGND VPWR VPWR _21334_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23216__A2 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24053_ _24488_/CLK _24053_/D HRESETn VGND VGND VPWR VPWR _13667_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21265_ _21275_/A _21263_/X _21265_/C VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__and3_4
X_23004_ _22801_/X _23002_/X _22804_/X _23003_/X VGND VGND VPWR VPWR _23005_/B sky130_fd_sc_hd__o22a_4
X_20216_ _20216_/A VGND VGND VPWR VPWR _20216_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21196_ _17714_/A _21194_/X _21195_/X VGND VGND VPWR VPWR _21196_/X sky130_fd_sc_hd__and3_4
XANTENNA__22090__A _22090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20147_ _20145_/Y _20141_/X _20146_/X _20129_/A VGND VGND VPWR VPWR _20147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_45_0_HCLK clkbuf_6_44_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20078_ _23524_/Q VGND VGND VPWR VPWR _20078_/Y sky130_fd_sc_hd__inv_2
X_24955_ _24979_/CLK _24955_/D HRESETn VGND VGND VPWR VPWR _24955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11920_ _11919_/X VGND VGND VPWR VPWR _11920_/Y sky130_fd_sc_hd__inv_2
X_23906_ _24214_/CLK _23906_/D VGND VGND VPWR VPWR _18985_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_218_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24886_ _24883_/CLK _24886_/D HRESETn VGND VGND VPWR VPWR _24886_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ _11851_/A VGND VGND VPWR VPWR _11851_/X sky130_fd_sc_hd__buf_2
XANTENNA__21434__A _22986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23837_ _23880_/CLK _23837_/D VGND VGND VPWR VPWR _19186_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_72_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19356__B1 _19220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11960__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _13575_/Y _14570_/B VGND VGND VPWR VPWR _14571_/B sky130_fd_sc_hd__or2_4
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _25547_/Q VGND VGND VPWR VPWR _11782_/Y sky130_fd_sc_hd__inv_2
X_23768_ _23768_/CLK _23768_/D VGND VGND VPWR VPWR _23768_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_HCLK clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _13516_/A VGND VGND VPWR VPWR _13521_/X sky130_fd_sc_hd__buf_2
X_25507_ _25507_/CLK _25507_/D HRESETn VGND VGND VPWR VPWR _25507_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_201_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22719_ _23253_/A _22719_/B _22718_/X VGND VGND VPWR VPWR _22719_/X sky130_fd_sc_hd__and3_4
XANTENNA__15917__B1 _15848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19839__A _19838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23699_ _23716_/CLK _23699_/D VGND VGND VPWR VPWR _23699_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ _13420_/A _23917_/Q VGND VGND VPWR VPWR _13454_/B sky130_fd_sc_hd__or2_4
X_16240_ _22716_/A VGND VGND VPWR VPWR _16240_/Y sky130_fd_sc_hd__inv_2
X_25438_ _25454_/CLK _25438_/D HRESETn VGND VGND VPWR VPWR _21083_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15932__A3 _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12403_/A VGND VGND VPWR VPWR _12403_/X sky130_fd_sc_hd__buf_2
X_13383_ _13310_/X _13381_/X _13382_/X VGND VGND VPWR VPWR _13383_/X sky130_fd_sc_hd__and3_4
X_16171_ _21531_/A VGND VGND VPWR VPWR _16171_/Y sky130_fd_sc_hd__inv_2
X_25369_ _25365_/CLK _13025_/X HRESETn VGND VGND VPWR VPWR _13023_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17359__A _17364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12334_ _25347_/Q _24832_/Q _12332_/Y _12333_/Y VGND VGND VPWR VPWR _12334_/X sky130_fd_sc_hd__o22a_4
X_15122_ _24990_/Q _15121_/A _15120_/Y _15121_/Y VGND VGND VPWR VPWR _15129_/B sky130_fd_sc_hd__o22a_4
XANTENNA__16342__B1 _16245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15053_ _14958_/Y VGND VGND VPWR VPWR _15053_/X sky130_fd_sc_hd__buf_2
X_19930_ _19930_/A VGND VGND VPWR VPWR _22094_/B sky130_fd_sc_hd__inv_2
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_255_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12265_ _12263_/Y _24757_/Q _25466_/Q _12264_/Y VGND VGND VPWR VPWR _12265_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22415__B1 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14004_ _14004_/A _14003_/Y VGND VGND VPWR VPWR _14004_/X sky130_fd_sc_hd__and2_4
XANTENNA__22712__B _22316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _19861_/A VGND VGND VPWR VPWR _19861_/Y sky130_fd_sc_hd__inv_2
X_12196_ _25454_/Q VGND VGND VPWR VPWR _12197_/A sky130_fd_sc_hd__inv_2
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18812_ _18630_/Y _18810_/X _18811_/Y VGND VGND VPWR VPWR _18812_/X sky130_fd_sc_hd__o21a_4
X_19792_ _23627_/Q VGND VGND VPWR VPWR _22233_/B sky130_fd_sc_hd__inv_2
XFILLER_96_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18743_ _18743_/A VGND VGND VPWR VPWR _18744_/B sky130_fd_sc_hd__inv_2
XFILLER_237_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15955_ _15938_/X _15943_/X HWDATA[26] _24779_/Q _15941_/X VGND VGND VPWR VPWR _15955_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14906_ _25029_/Q VGND VGND VPWR VPWR _14906_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18674_ _18652_/X _18659_/X _18667_/X _18673_/X VGND VGND VPWR VPWR _18674_/X sky130_fd_sc_hd__or4_4
X_15886_ _12833_/Y _15880_/X _11783_/X _15880_/X VGND VGND VPWR VPWR _15886_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17625_ _17573_/A _17627_/B _17624_/Y VGND VGND VPWR VPWR _24321_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21344__A _23148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14837_ _14837_/A VGND VGND VPWR VPWR _14837_/X sky130_fd_sc_hd__buf_2
XANTENNA__25308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11870__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17556_ _11859_/Y _24299_/Q _11869_/A _17537_/Y VGND VGND VPWR VPWR _17560_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_65_0_HCLK clkbuf_7_32_0_HCLK/X VGND VGND VPWR VPWR _25454_/CLK sky130_fd_sc_hd__clkbuf_1
X_14768_ _21629_/A _14755_/B _14761_/X VGND VGND VPWR VPWR _25066_/D sky130_fd_sc_hd__a21oi_4
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21154__B1 _21583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16507_ _16540_/A VGND VGND VPWR VPWR _16533_/A sky130_fd_sc_hd__buf_2
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13719_ _11688_/Y _13699_/B VGND VGND VPWR VPWR _13719_/Y sky130_fd_sc_hd__nand2_4
X_17487_ _17486_/X VGND VGND VPWR VPWR _17487_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14699_ _13757_/A _14761_/A _13757_/A _14761_/A VGND VGND VPWR VPWR _14728_/A sky130_fd_sc_hd__a2bb2o_4
X_19226_ _19091_/A VGND VGND VPWR VPWR _19226_/X sky130_fd_sc_hd__buf_2
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16438_ _16442_/A VGND VGND VPWR VPWR _16438_/X sky130_fd_sc_hd__buf_2
XFILLER_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22675__A1_N _22678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19157_ _19156_/Y _19152_/X _19131_/X _19152_/X VGND VGND VPWR VPWR _23848_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17269__A _17345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16369_ _16367_/Y _16365_/X _16368_/X _16365_/X VGND VGND VPWR VPWR _16369_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18108_ _15704_/X _18088_/X _18107_/X _24252_/Q _18029_/X VGND VGND VPWR VPWR _18108_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__24943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19088_ _19087_/Y _19082_/X _18991_/X _19082_/X VGND VGND VPWR VPWR _19088_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18039_ _18039_/A _19330_/A VGND VGND VPWR VPWR _18039_/X sky130_fd_sc_hd__or2_4
XFILLER_172_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16901__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21050_ _21024_/B _21105_/B VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__and2_4
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21519__A _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22421__A3 _21308_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20001_ _21956_/B _19997_/X _20000_/X _19997_/X VGND VGND VPWR VPWR _20001_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21952_ _21473_/A _21952_/B VGND VGND VPWR VPWR _21952_/X sky130_fd_sc_hd__or2_4
X_24740_ _24738_/CLK _16037_/X HRESETn VGND VGND VPWR VPWR _24740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_228_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20903_ _24062_/Q _20897_/X _20911_/B VGND VGND VPWR VPWR _20903_/Y sky130_fd_sc_hd__a21oi_4
X_24671_ _24552_/CLK _16228_/X HRESETn VGND VGND VPWR VPWR _16226_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_242_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21883_ _24794_/Q _21881_/X _22954_/C _24864_/Q _21085_/A VGND VGND VPWR VPWR _21883_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_215_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16348__A _16348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11780__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23622_ _23597_/CLK _23622_/D VGND VGND VPWR VPWR _23622_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_243_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20834_ _20831_/A _20834_/B VGND VGND VPWR VPWR _20842_/A sky130_fd_sc_hd__or2_4
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21145__B1 _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _23553_/CLK _20001_/X VGND VGND VPWR VPWR _23553_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20765_ _20765_/A VGND VGND VPWR VPWR _20765_/X sky130_fd_sc_hd__buf_2
XANTENNA__19659__A _19151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _15800_/A _22502_/X _22503_/X _25534_/Q _16003_/A VGND VGND VPWR VPWR _22504_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _23516_/CLK _20194_/X VGND VGND VPWR VPWR _20190_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20696_ _20693_/A _20696_/B VGND VGND VPWR VPWR _20724_/A sky130_fd_sc_hd__or2_4
XFILLER_149_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15914__A3 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25223_ _25223_/CLK _25223_/D HRESETn VGND VGND VPWR VPWR _14110_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_155_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22435_ _22401_/X _22435_/B _22435_/C _22435_/D VGND VGND VPWR VPWR HRDATA[7] sky130_fd_sc_hd__or4_4
XANTENNA__22645__B1 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24684__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25154_ _25154_/CLK _25154_/D HRESETn VGND VGND VPWR VPWR _25154_/Q sky130_fd_sc_hd__dfrtp_4
X_22366_ _21948_/A _22366_/B VGND VGND VPWR VPWR _22366_/X sky130_fd_sc_hd__or2_4
XFILLER_108_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20120__B2 _20118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24105_ _23631_/CLK _20973_/X HRESETn VGND VGND VPWR VPWR _24105_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24613__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21317_ _21316_/X VGND VGND VPWR VPWR _21317_/X sky130_fd_sc_hd__buf_2
X_25085_ _25062_/CLK _25085_/D HRESETn VGND VGND VPWR VPWR _14624_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22297_ _16713_/Y _22424_/B VGND VGND VPWR VPWR _22297_/X sky130_fd_sc_hd__and2_4
XANTENNA__16811__A _16810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12050_ _12050_/A VGND VGND VPWR VPWR _12050_/X sky130_fd_sc_hd__buf_2
X_24036_ _24500_/CLK _20793_/X HRESETn VGND VGND VPWR VPWR _20789_/A sky130_fd_sc_hd__dfrtp_4
X_21248_ _21248_/A VGND VGND VPWR VPWR _21271_/A sky130_fd_sc_hd__buf_2
XANTENNA__21429__A _21535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19813__B2 _19788_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11955__A _19643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21179_ _17455_/X VGND VGND VPWR VPWR _22527_/A sky130_fd_sc_hd__inv_2
XFILLER_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15740_ _12595_/Y _15730_/X _11783_/X _15730_/X VGND VGND VPWR VPWR _15740_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15850__A2 _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12952_ _12783_/Y _12969_/A _12952_/C _12952_/D VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__or4_4
X_24938_ _24937_/CLK _24938_/D HRESETn VGND VGND VPWR VPWR _11740_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_234_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20187__B2 _20184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22581__C1 _22580_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11903_ _11933_/A _11898_/A VGND VGND VPWR VPWR _11903_/X sky130_fd_sc_hd__and2_4
X_15671_ _21140_/A _17448_/C _21045_/A _15670_/X VGND VGND VPWR VPWR _21170_/A sky130_fd_sc_hd__or4_4
XANTENNA__11872__B1 _11871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12883_ _12908_/A VGND VGND VPWR VPWR _12883_/X sky130_fd_sc_hd__buf_2
X_24869_ _24867_/CLK _24869_/D HRESETn VGND VGND VPWR VPWR _24869_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19329__B1 _19305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17410_/A VGND VGND VPWR VPWR _17410_/X sky130_fd_sc_hd__buf_2
XPHY_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _25086_/Q VGND VGND VPWR VPWR _14622_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11834_ HWDATA[9] VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__buf_2
X_18390_ _24198_/Q VGND VGND VPWR VPWR _18390_/Y sky130_fd_sc_hd__inv_2
XPHY_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A _17341_/B VGND VGND VPWR VPWR _17342_/C sky130_fd_sc_hd__or2_4
XFILLER_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _25552_/Q VGND VGND VPWR VPWR _11765_/Y sky130_fd_sc_hd__inv_2
X_14553_ _14553_/A VGND VGND VPWR VPWR _14554_/C sky130_fd_sc_hd__inv_2
XANTENNA__22884__B1 _25543_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22707__B _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _16193_/A _13504_/B VGND VGND VPWR VPWR _13504_/X sky130_fd_sc_hd__or2_4
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _24377_/Q _17271_/Y VGND VGND VPWR VPWR _17272_/X sky130_fd_sc_hd__or2_4
XFILLER_158_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11694_/A _24239_/Q _13697_/A _11695_/Y VGND VGND VPWR VPWR _11697_/D sky130_fd_sc_hd__o22a_4
X_14484_ _14484_/A _14416_/X VGND VGND VPWR VPWR _14485_/A sky130_fd_sc_hd__nor2_4
XANTENNA__16563__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ HWDATA[5] VGND VGND VPWR VPWR _19151_/A sky130_fd_sc_hd__buf_2
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16223_ _16221_/Y _16222_/X _15963_/X _16222_/X VGND VGND VPWR VPWR _16223_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13435_ _13371_/A _13435_/B VGND VGND VPWR VPWR _13435_/X sky130_fd_sc_hd__or2_4
XFILLER_173_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12952__C _12952_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13290_/X _13366_/B _13365_/X VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__and3_4
X_16154_ _16162_/A VGND VGND VPWR VPWR _16154_/X sky130_fd_sc_hd__buf_2
XFILLER_10_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _24604_/Q VGND VGND VPWR VPWR _15105_/Y sky130_fd_sc_hd__inv_2
X_12317_ _12317_/A VGND VGND VPWR VPWR _12317_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13297_ _13369_/A _13297_/B VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__or2_4
X_16085_ _16084_/Y _16005_/X _15489_/X _16005_/X VGND VGND VPWR VPWR _16085_/X sky130_fd_sc_hd__a2bb2o_4
X_12248_ _12247_/X _24767_/Q _12247_/A _24767_/Q VGND VGND VPWR VPWR _12249_/D sky130_fd_sc_hd__a2bb2o_4
X_15036_ _15036_/A VGND VGND VPWR VPWR _15036_/Y sky130_fd_sc_hd__inv_2
X_19913_ _21955_/B _19910_/X _19636_/X _19910_/X VGND VGND VPWR VPWR _23585_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20243__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12352__B2 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11865__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19844_ _19838_/Y VGND VGND VPWR VPWR _19844_/X sky130_fd_sc_hd__buf_2
X_12179_ _12168_/X _12178_/X SCLK_S3 _12168_/X VGND VGND VPWR VPWR _12179_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19775_ _23633_/Q VGND VGND VPWR VPWR _19775_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15056__B _15052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16784__A1_N _15017_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ _24385_/Q VGND VGND VPWR VPWR _16987_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18726_ _24158_/Q _18725_/Y VGND VGND VPWR VPWR _18726_/X sky130_fd_sc_hd__or2_4
X_15938_ _15796_/X VGND VGND VPWR VPWR _15938_/X sky130_fd_sc_hd__buf_2
XANTENNA__20178__B2 _20177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18657_ _24146_/Q VGND VGND VPWR VPWR _18657_/X sky130_fd_sc_hd__buf_2
XANTENNA__11863__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15869_ _21069_/B VGND VGND VPWR VPWR _15870_/B sky130_fd_sc_hd__buf_2
X_17608_ _17598_/A _17608_/B _17607_/X VGND VGND VPWR VPWR _17608_/X sky130_fd_sc_hd__and3_4
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18588_ _18434_/A _18588_/B VGND VGND VPWR VPWR _18588_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_10_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17539_ _11869_/A _17537_/Y _25530_/Q _17588_/A VGND VGND VPWR VPWR _17542_/B sky130_fd_sc_hd__a2bb2o_4
X_20550_ _18891_/X VGND VGND VPWR VPWR _20550_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_9_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19209_ _17951_/B VGND VGND VPWR VPWR _19209_/Y sky130_fd_sc_hd__inv_2
X_20481_ _20609_/B _20480_/X _14550_/A _20443_/X VGND VGND VPWR VPWR _24094_/D sky130_fd_sc_hd__a211o_4
XFILLER_165_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22220_ _22209_/A _22218_/X _22220_/C VGND VGND VPWR VPWR _22220_/X sky130_fd_sc_hd__and3_4
XANTENNA__13320__A _13320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15109__B2 _15108_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18846__A2 _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22642__A3 _22303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22151_ _21872_/A VGND VGND VPWR VPWR _23093_/A sky130_fd_sc_hd__buf_2
XANTENNA__21850__A1 _20525_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21102_ _15866_/X VGND VGND VPWR VPWR _21103_/A sky130_fd_sc_hd__buf_2
X_22082_ _22394_/A _20133_/Y VGND VGND VPWR VPWR _22083_/C sky130_fd_sc_hd__or2_4
XFILLER_161_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_221_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21033_ _21032_/X VGND VGND VPWR VPWR _21605_/A sky130_fd_sc_hd__buf_2
XFILLER_160_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13540__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22158__A2 _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22984_ _23117_/A _22983_/X VGND VGND VPWR VPWR _22984_/X sky130_fd_sc_hd__and2_4
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24723_ _24735_/CLK _16081_/X HRESETn VGND VGND VPWR VPWR _24723_/Q sky130_fd_sc_hd__dfrtp_4
X_21935_ _21209_/A VGND VGND VPWR VPWR _21945_/A sky130_fd_sc_hd__buf_2
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21866_ _21584_/X _21864_/X _21578_/X _21865_/X VGND VGND VPWR VPWR _21866_/X sky130_fd_sc_hd__o22a_4
X_24654_ _24194_/CLK _24654_/D HRESETn VGND VGND VPWR VPWR _16273_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_203_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16793__B1 _16791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20822_/B VGND VGND VPWR VPWR _20818_/A sky130_fd_sc_hd__inv_2
X_23605_ _23597_/CLK _23605_/D VGND VGND VPWR VPWR _23605_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21712__A _21712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21654_/X _21796_/X _25279_/Q _18268_/X VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__o22a_4
X_24585_ _24556_/CLK _16455_/X HRESETn VGND VGND VPWR VPWR _24585_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19731__B1 _19612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24865__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15710__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20748_ _20739_/X _20747_/X _15618_/A _20744_/X VGND VGND VPWR VPWR _20748_/X sky130_fd_sc_hd__a2bb2o_4
X_23536_ _23560_/CLK _23536_/D VGND VGND VPWR VPWR _23536_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16545__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20341__B2 _20323_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23794_/CLK _23467_/D VGND VGND VPWR VPWR _17987_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_195_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20679_ _14227_/Y _17413_/A _17396_/A _17410_/A VGND VGND VPWR VPWR _20679_/X sky130_fd_sc_hd__o22a_4
XFILLER_109_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13420_/A _13220_/B VGND VGND VPWR VPWR _13220_/X sky130_fd_sc_hd__or2_4
X_22418_ _22418_/A _22284_/X VGND VGND VPWR VPWR _22418_/X sky130_fd_sc_hd__or2_4
X_25206_ _24000_/CLK _14234_/X HRESETn VGND VGND VPWR VPWR _14227_/A sky130_fd_sc_hd__dfstp_4
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23398_ _24206_/CLK _23398_/D VGND VGND VPWR VPWR _23398_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22543__A _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13151_ _21130_/A _13149_/X _13150_/Y VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__o21a_4
X_22349_ _22345_/X _22348_/X _17732_/A VGND VGND VPWR VPWR _22349_/Y sky130_fd_sc_hd__o21ai_4
X_25137_ _25137_/CLK _25137_/D HRESETn VGND VGND VPWR VPWR _25137_/Q sky130_fd_sc_hd__dfstp_4
X_12102_ _13798_/B VGND VGND VPWR VPWR _12102_/X sky130_fd_sc_hd__buf_2
X_13082_ _13084_/B VGND VGND VPWR VPWR _13083_/B sky130_fd_sc_hd__inv_2
X_25068_ _25068_/CLK _25068_/D HRESETn VGND VGND VPWR VPWR _25068_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23043__B1 _12595_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12033_ _24109_/Q _12024_/X _12030_/Y VGND VGND VPWR VPWR _20977_/A sky130_fd_sc_hd__o21a_4
X_16910_ _16910_/A VGND VGND VPWR VPWR _16910_/Y sky130_fd_sc_hd__inv_2
X_24019_ _24020_/CLK _20715_/Y HRESETn VGND VGND VPWR VPWR _13135_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_239_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17890_ _17758_/Y _17888_/X _17889_/Y VGND VGND VPWR VPWR _17890_/X sky130_fd_sc_hd__o21a_4
X_16841_ _16841_/A VGND VGND VPWR VPWR _16841_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23374__A _23361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15284__B1 _14996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19560_ _11855_/A VGND VGND VPWR VPWR _19560_/X sky130_fd_sc_hd__buf_2
XFILLER_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12098__B1 _11871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16772_ _22713_/A VGND VGND VPWR VPWR _16772_/Y sky130_fd_sc_hd__inv_2
X_13984_ _13984_/A VGND VGND VPWR VPWR _14058_/A sky130_fd_sc_hd__buf_2
X_18511_ _18492_/A _18509_/X _18510_/X VGND VGND VPWR VPWR _18511_/X sky130_fd_sc_hd__and3_4
X_15723_ HWDATA[30] VGND VGND VPWR VPWR _15723_/X sky130_fd_sc_hd__buf_2
X_12935_ _25388_/Q _12934_/Y VGND VGND VPWR VPWR _12935_/X sky130_fd_sc_hd__or2_4
X_19491_ _19491_/A VGND VGND VPWR VPWR _21959_/B sky130_fd_sc_hd__inv_2
XFILLER_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18442_ _16237_/Y _24178_/Q _16237_/Y _24178_/Q VGND VGND VPWR VPWR _18443_/D sky130_fd_sc_hd__a2bb2o_4
X_15654_ _15657_/A VGND VGND VPWR VPWR _21299_/A sky130_fd_sc_hd__inv_2
XFILLER_61_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12866_ _12790_/Y _12878_/A _12839_/Y _12865_/X VGND VGND VPWR VPWR _12869_/B sky130_fd_sc_hd__or4_4
XANTENNA__16784__B1 _16613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14605_ _14605_/A _14574_/X VGND VGND VPWR VPWR _14605_/Y sky130_fd_sc_hd__nand2_4
XPHY_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ HWDATA[13] VGND VGND VPWR VPWR _16245_/A sky130_fd_sc_hd__buf_2
X_18373_ _18361_/X _18359_/Y _18372_/X _18357_/A _18362_/Y VGND VGND VPWR VPWR _24205_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15583_/Y _15584_/X _11773_/X _15584_/X VGND VGND VPWR VPWR _15585_/X sky130_fd_sc_hd__a2bb2o_4
X_12797_ _21537_/A VGND VGND VPWR VPWR _12797_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17229_/Y _17318_/X _17288_/X _17321_/B VGND VGND VPWR VPWR _17324_/X sky130_fd_sc_hd__a211o_4
X_14536_ _14530_/X _14535_/X _14494_/A _14526_/X VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__o22a_4
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11730_/Y _22694_/B VGND VGND VPWR VPWR _11749_/A sky130_fd_sc_hd__and2_4
XFILLER_187_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_139_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _25082_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _17205_/Y _17193_/Y _17184_/A _17255_/D VGND VGND VPWR VPWR _17256_/D sky130_fd_sc_hd__or4_4
XFILLER_174_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22609__B1 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14467_ _14467_/A VGND VGND VPWR VPWR _14467_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11679_ _13736_/A _24234_/Q _13736_/A _24234_/Q VGND VGND VPWR VPWR _11684_/B sky130_fd_sc_hd__a2bb2o_4
X_16206_ _16205_/Y _16203_/X _15950_/X _16203_/X VGND VGND VPWR VPWR _16206_/X sky130_fd_sc_hd__a2bb2o_4
X_13418_ _13450_/A _23910_/Q VGND VGND VPWR VPWR _13419_/C sky130_fd_sc_hd__or2_4
X_17186_ _17186_/A VGND VGND VPWR VPWR _17322_/A sky130_fd_sc_hd__inv_2
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23282__B1 _11757_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14398_ _20470_/A _14391_/X _13849_/X _14393_/X VGND VGND VPWR VPWR _14398_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20096__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16137_ _16134_/Y _16136_/X _11805_/X _16136_/X VGND VGND VPWR VPWR _24702_/D sky130_fd_sc_hd__a2bb2o_4
X_13349_ _13413_/A _13349_/B VGND VGND VPWR VPWR _13349_/X sky130_fd_sc_hd__or2_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16451__A _19091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22172__B _22316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16068_ _24727_/Q VGND VGND VPWR VPWR _16068_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13522__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15019_ _15019_/A VGND VGND VPWR VPWR _15019_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19827_ _19826_/Y _19822_/X _19753_/X _19822_/X VGND VGND VPWR VPWR _23616_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23337__A1 _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18378__A _18377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12089__B1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19758_ _13433_/B VGND VGND VPWR VPWR _19758_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18709_ _18739_/A _18709_/B _18709_/C VGND VGND VPWR VPWR _18709_/X sky130_fd_sc_hd__and3_4
XANTENNA__11836__B1 _11834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19689_ _19675_/Y VGND VGND VPWR VPWR _19689_/X sky130_fd_sc_hd__buf_2
XFILLER_225_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21720_ _22289_/A _21719_/X _21550_/X _16078_/A _21551_/X VGND VGND VPWR VPWR _21720_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13315__A _13315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22560__A2 _23303_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19961__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16775__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21651_ _14725_/X _21651_/B _21650_/X VGND VGND VPWR VPWR _21651_/X sky130_fd_sc_hd__or3_4
XFILLER_224_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_35_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_70_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20602_ _18887_/A _18887_/B _20601_/Y _20550_/Y VGND VGND VPWR VPWR _20603_/C sky130_fd_sc_hd__a211o_4
X_24370_ _24372_/CLK _24370_/D HRESETn VGND VGND VPWR VPWR _17195_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_33_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21582_ _18390_/Y _21580_/X _12127_/Y _21579_/X VGND VGND VPWR VPWR _21582_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_98_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_98_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22863__A3 _22861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23321_ _23321_/A _23320_/X VGND VGND VPWR VPWR _23331_/B sky130_fd_sc_hd__and2_4
XFILLER_193_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20533_ _23979_/Q _14290_/A _20533_/C _20532_/X VGND VGND VPWR VPWR _20534_/A sky130_fd_sc_hd__or4_4
XFILLER_178_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23252_ _16562_/A _22485_/X _22852_/X _23251_/X VGND VGND VPWR VPWR _23253_/C sky130_fd_sc_hd__a211o_4
X_20464_ _20462_/X _20463_/X VGND VGND VPWR VPWR _20464_/X sky130_fd_sc_hd__or2_4
XFILLER_229_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22203_ _25531_/Q _22425_/B _21121_/A _22202_/X VGND VGND VPWR VPWR _22204_/C sky130_fd_sc_hd__a211o_4
XANTENNA__20087__B1 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23183_ _23183_/A _23183_/B VGND VGND VPWR VPWR _23187_/B sky130_fd_sc_hd__or2_4
XFILLER_180_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17457__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20395_ _23407_/Q VGND VGND VPWR VPWR _21818_/B sky130_fd_sc_hd__inv_2
XANTENNA__16361__A _24622_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_HCLK clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21575__A2_N _16192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22134_ _20525_/A _22176_/B _23974_/Q _21369_/B VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13513__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12316__B2 _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22065_ _19556_/Y _22013_/Y _22014_/X _22064_/X VGND VGND VPWR VPWR _22066_/A sky130_fd_sc_hd__a211o_4
XFILLER_181_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21016_ _21016_/A VGND VGND VPWR VPWR _21018_/B sky130_fd_sc_hd__inv_2
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15266__B1 _14996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18288__A _17712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16614__A1_N _16612_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22967_ _24605_/Q _22849_/X VGND VGND VPWR VPWR _22967_/X sky130_fd_sc_hd__or2_4
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _12623_/C _12722_/B _12719_/Y VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__o21a_4
X_24706_ _24712_/CLK _24706_/D HRESETn VGND VGND VPWR VPWR _24706_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13225__A _13315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21918_ _21895_/X _20200_/Y VGND VGND VPWR VPWR _21918_/X sky130_fd_sc_hd__or2_4
XANTENNA__16766__B1 _16419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22898_ _24570_/Q _22897_/X _22816_/X VGND VGND VPWR VPWR _22898_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21442__A _15866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12651_ _12702_/A _12642_/D VGND VGND VPWR VPWR _12654_/B sky130_fd_sc_hd__or2_4
X_24637_ _24629_/CLK _24637_/D HRESETn VGND VGND VPWR VPWR _16322_/A sky130_fd_sc_hd__dfrtp_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21849_ _14240_/Y _14232_/A _15479_/Y _15471_/A VGND VGND VPWR VPWR _21851_/B sky130_fd_sc_hd__o22a_4
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__A _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12660_/A _24883_/Q _12660_/A _24883_/Q VGND VGND VPWR VPWR _12582_/X sky130_fd_sc_hd__a2bb2o_4
X_15370_ _15370_/A _15369_/X VGND VGND VPWR VPWR _15384_/B sky130_fd_sc_hd__or2_4
XANTENNA__16518__B1 _16248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12252__B1 _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24568_ _24592_/CLK _16509_/X HRESETn VGND VGND VPWR VPWR _16506_/A sky130_fd_sc_hd__dfrtp_4
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _14315_/X _14319_/X _25328_/Q _14320_/X VGND VGND VPWR VPWR _14321_/X sky130_fd_sc_hd__o22a_4
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23519_ _23918_/CLK _20094_/X VGND VGND VPWR VPWR _23519_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24499_ _24532_/CLK _16693_/X HRESETn VGND VGND VPWR VPWR _24499_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _24393_/Q VGND VGND VPWR VPWR _17042_/C sky130_fd_sc_hd__inv_2
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22067__A1 _25265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _13924_/D VGND VGND VPWR VPWR _14252_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22606__A3 _22145_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13203_ _11973_/A _11984_/C VGND VGND VPWR VPWR _13203_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17367__A _17364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14183_ _14179_/Y _14182_/Y _14174_/X VGND VGND VPWR VPWR _14183_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ _24018_/Q _13134_/B VGND VGND VPWR VPWR _13134_/X sky130_fd_sc_hd__or2_4
X_18991_ _19131_/A VGND VGND VPWR VPWR _18991_/X sky130_fd_sc_hd__buf_2
XANTENNA__12307__B2 _24852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13065_ _12323_/Y _13069_/B _13064_/Y VGND VGND VPWR VPWR _25359_/D sky130_fd_sc_hd__o21a_4
X_17942_ _18023_/A VGND VGND VPWR VPWR _17943_/A sky130_fd_sc_hd__buf_2
XFILLER_78_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22720__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12016_ _13514_/A _12015_/Y _13514_/A _12015_/Y VGND VGND VPWR VPWR _12021_/C sky130_fd_sc_hd__a2bb2o_4
X_17873_ _17881_/A _17873_/B _17873_/C VGND VGND VPWR VPWR _24272_/D sky130_fd_sc_hd__and3_4
XFILLER_94_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20250__B1 _20249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16824_ _14980_/Y _16820_/X HWDATA[22] _16820_/X VGND VGND VPWR VPWR _16824_/X sky130_fd_sc_hd__a2bb2o_4
X_19612_ _11861_/A VGND VGND VPWR VPWR _19612_/X sky130_fd_sc_hd__buf_2
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19543_ _23710_/Q VGND VGND VPWR VPWR _21502_/B sky130_fd_sc_hd__inv_2
X_16755_ _16754_/Y _16752_/X _15738_/X _16752_/X VGND VGND VPWR VPWR _16755_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _13967_/A _13967_/B _13967_/C _13899_/X VGND VGND VPWR VPWR _13967_/X sky130_fd_sc_hd__or4_4
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15706_ _24893_/Q _15700_/Y _15696_/C _15705_/X VGND VGND VPWR VPWR _15706_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24787__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12918_ _12927_/A _12916_/X _12918_/C VGND VGND VPWR VPWR _25394_/D sky130_fd_sc_hd__and3_4
X_19474_ _19472_/Y _19473_/X _19383_/X _19473_/X VGND VGND VPWR VPWR _23735_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16686_ _16684_/Y _16680_/X _16417_/X _16685_/X VGND VGND VPWR VPWR _24502_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16757__B1 _16407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20553__A1 _14178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13898_ _13928_/A _13929_/A _13950_/A _13952_/C VGND VGND VPWR VPWR _13899_/C sky130_fd_sc_hd__or4_4
XFILLER_179_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18425_ _24165_/Q VGND VGND VPWR VPWR _18425_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24716__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _15634_/Y _15635_/X _15636_/X _15635_/X VGND VGND VPWR VPWR _24903_/D sky130_fd_sc_hd__a2bb2o_4
X_12849_ _25401_/Q VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__inv_2
XANTENNA__16446__A _16390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22167__B _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_2_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _18355_/Y _18361_/A _24206_/Q _17492_/X VGND VGND VPWR VPWR _18370_/A sky130_fd_sc_hd__o22a_4
XFILLER_194_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15568_ _24928_/Q VGND VGND VPWR VPWR _15568_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16509__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17307_ _17248_/B _17301_/X _17288_/X _17303_/Y VGND VGND VPWR VPWR _17308_/A sky130_fd_sc_hd__a211o_4
X_14519_ _23970_/Q VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__buf_2
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18287_ _18286_/Y VGND VGND VPWR VPWR _20015_/B sky130_fd_sc_hd__buf_2
XFILLER_174_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15499_ _15499_/A VGND VGND VPWR VPWR _15503_/A sky130_fd_sc_hd__buf_2
XFILLER_175_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17238_ _17238_/A _17235_/X _17236_/X _17238_/D VGND VGND VPWR VPWR _17239_/D sky130_fd_sc_hd__or4_4
XFILLER_174_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17169_ _17166_/B _17168_/Y _17160_/C VGND VGND VPWR VPWR _17169_/X sky130_fd_sc_hd__and3_4
X_20180_ _20179_/Y _20177_/X _20112_/X _20177_/X VGND VGND VPWR VPWR _23489_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21569__B1 _14877_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20241__B1 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23870_ _23871_/CLK _19094_/X VGND VGND VPWR VPWR _23870_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22821_ _16506_/A _22543_/A _22544_/X VGND VGND VPWR VPWR _22821_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25540_ _25539_/CLK _25540_/D HRESETn VGND VGND VPWR VPWR _25540_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22752_ _16510_/A _22543_/X _22545_/X VGND VGND VPWR VPWR _22752_/X sky130_fd_sc_hd__o21a_4
XFILLER_198_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21703_ _21513_/X _21702_/X _11703_/Y _21513_/X VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22683_ _16841_/Y _21431_/X _21591_/X _22682_/X VGND VGND VPWR VPWR _22683_/X sky130_fd_sc_hd__o22a_4
X_25471_ _24196_/CLK _12183_/X HRESETn VGND VGND VPWR VPWR _25471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16356__A _24624_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21634_ _22388_/A _20183_/Y VGND VGND VPWR VPWR _21637_/B sky130_fd_sc_hd__or2_4
X_24422_ _24613_/CLK _24422_/D HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_240_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12785__A1 _25380_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21565_ _21565_/A VGND VGND VPWR VPWR _21565_/Y sky130_fd_sc_hd__inv_2
X_24353_ _24354_/CLK _17377_/X HRESETn VGND VGND VPWR VPWR _24353_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19667__A _19652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22805__B _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20516_ _24013_/Q _20456_/X _20515_/X VGND VGND VPWR VPWR _24013_/D sky130_fd_sc_hd__a21o_4
X_23304_ _15568_/Y _22890_/B VGND VGND VPWR VPWR _23304_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_122_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24500_/CLK sky130_fd_sc_hd__clkbuf_1
X_24284_ _24283_/CLK _17825_/X HRESETn VGND VGND VPWR VPWR _16909_/A sky130_fd_sc_hd__dfrtp_4
X_21496_ _22271_/A VGND VGND VPWR VPWR _21497_/A sky130_fd_sc_hd__buf_2
XANTENNA__22093__A _22093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_185_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _25168_/CLK sky130_fd_sc_hd__clkbuf_1
X_23235_ _23124_/X _23234_/X _23058_/X _24749_/Q _21538_/X VGND VGND VPWR VPWR _23236_/A
+ sky130_fd_sc_hd__a32o_4
X_20447_ _20446_/X VGND VGND VPWR VPWR _20447_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23166_ _23124_/X _23165_/X _23058_/X _16018_/A _22990_/X VGND VGND VPWR VPWR _23167_/A
+ sky130_fd_sc_hd__a32o_4
X_20378_ _21672_/B _20377_/X _19643_/A _20377_/X VGND VGND VPWR VPWR _20378_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15487__B1 _15486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22117_ _22117_/A VGND VGND VPWR VPWR _22119_/C sky130_fd_sc_hd__inv_2
X_23097_ _16669_/Y _22842_/X _15586_/Y _22845_/X VGND VGND VPWR VPWR _23097_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22540__B _22589_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22048_ _21682_/A _19909_/Y _21685_/X VGND VGND VPWR VPWR _22048_/X sky130_fd_sc_hd__o21a_4
XFILLER_76_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12252__A1_N _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21437__A _21436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22772__A2 _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14870_ _14822_/C _14822_/B _14822_/C _14822_/B VGND VGND VPWR VPWR _14870_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13821_ _17448_/A _13821_/B VGND VGND VPWR VPWR _13822_/B sky130_fd_sc_hd__or2_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23999_ _25246_/CLK _20678_/Y HRESETn VGND VGND VPWR VPWR _23999_/Q sky130_fd_sc_hd__dfrtp_4
X_16540_ _16540_/A VGND VGND VPWR VPWR _16540_/X sky130_fd_sc_hd__buf_2
XFILLER_244_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17650__A _17578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24880__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13752_ _13749_/Y _13751_/Y VGND VGND VPWR VPWR _14789_/A sky130_fd_sc_hd__or2_4
XFILLER_232_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _12574_/Y _12702_/X VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__or2_4
XFILLER_243_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21172__A _16864_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16471_ _16466_/Y _16470_/X _16385_/X _16470_/X VGND VGND VPWR VPWR _24583_/D sky130_fd_sc_hd__a2bb2o_4
X_13683_ _25303_/Q _13533_/X _13682_/Y VGND VGND VPWR VPWR _13683_/X sky130_fd_sc_hd__o21a_4
X_18210_ _18178_/A _20253_/A VGND VGND VPWR VPWR _18211_/C sky130_fd_sc_hd__or2_4
XFILLER_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15422_ _15421_/X VGND VGND VPWR VPWR _15422_/Y sky130_fd_sc_hd__inv_2
X_12634_ _12521_/A _12633_/Y VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__or2_4
X_19190_ _19189_/X VGND VGND VPWR VPWR _19196_/A sky130_fd_sc_hd__inv_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18141_ _17973_/X _18140_/X _24250_/Q _18031_/X VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12820__A1_N _12819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15353_ _15346_/B VGND VGND VPWR VPWR _15357_/B sky130_fd_sc_hd__inv_2
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12563_/A _24878_/Q _12619_/A _12564_/Y VGND VGND VPWR VPWR _12565_/X sky130_fd_sc_hd__o22a_4
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_81_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _14304_/A VGND VGND VPWR VPWR _14316_/A sky130_fd_sc_hd__buf_2
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18072_ _13613_/B VGND VGND VPWR VPWR _18072_/X sky130_fd_sc_hd__buf_2
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _15258_/A _15257_/X _14996_/X _15282_/B VGND VGND VPWR VPWR _15285_/A sky130_fd_sc_hd__a211o_4
XFILLER_184_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12238_/Y _12502_/A VGND VGND VPWR VPWR _12500_/B sky130_fd_sc_hd__or2_4
X_17023_ _24749_/Q _17034_/A _16075_/Y _17051_/A VGND VGND VPWR VPWR _17025_/C sky130_fd_sc_hd__a2bb2o_4
X_14235_ _25205_/Q VGND VGND VPWR VPWR _14235_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17097__A _17393_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14166_ _14138_/X _14165_/X _25141_/Q _14145_/X VGND VGND VPWR VPWR _14166_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__18664__B1 _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15478__B1 _14427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13117_ _12387_/X _13121_/A VGND VGND VPWR VPWR _13117_/Y sky130_fd_sc_hd__nand2_4
X_14097_ _13994_/B _14090_/X _14078_/X _13994_/A _14093_/X VGND VGND VPWR VPWR _14097_/X
+ sky130_fd_sc_hd__a32o_4
X_18974_ _18974_/A VGND VGND VPWR VPWR _18974_/X sky130_fd_sc_hd__buf_2
XFILLER_79_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13048_ _13007_/X _13026_/D _12370_/Y VGND VGND VPWR VPWR _13049_/C sky130_fd_sc_hd__o21a_4
X_17925_ _13550_/X VGND VGND VPWR VPWR _17925_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23265__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15345__A _15388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11873__A _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17856_ _16916_/Y VGND VGND VPWR VPWR _17861_/B sky130_fd_sc_hd__buf_2
XANTENNA__21066__B _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17263__C _17263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16807_ _16803_/Y _16806_/X _16385_/X _16806_/X VGND VGND VPWR VPWR _24450_/D sky130_fd_sc_hd__a2bb2o_4
X_17787_ _17787_/A _17787_/B VGND VGND VPWR VPWR _17789_/B sky130_fd_sc_hd__or2_4
XFILLER_226_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14999_ _25014_/Q VGND VGND VPWR VPWR _15292_/A sky130_fd_sc_hd__inv_2
XFILLER_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16738_ _16737_/Y VGND VGND VPWR VPWR _16738_/X sky130_fd_sc_hd__buf_2
X_19526_ _23716_/Q VGND VGND VPWR VPWR _22358_/B sky130_fd_sc_hd__inv_2
XANTENNA__21723__B1 _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24550__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19457_ _19456_/Y _19451_/X _19410_/X _19438_/A VGND VGND VPWR VPWR _23741_/D sky130_fd_sc_hd__a2bb2o_4
X_16669_ _16669_/A VGND VGND VPWR VPWR _16669_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18408_ _24190_/Q VGND VGND VPWR VPWR _18510_/A sky130_fd_sc_hd__inv_2
X_19388_ _19387_/Y _19382_/X _19254_/X _19368_/Y VGND VGND VPWR VPWR _23765_/D sky130_fd_sc_hd__a2bb2o_4
X_18339_ _18937_/B VGND VGND VPWR VPWR _20079_/C sky130_fd_sc_hd__buf_2
XANTENNA__25147__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12209__A _22871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21350_ _21731_/A VGND VGND VPWR VPWR _21350_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20301_ _19965_/A _19986_/X _18289_/X VGND VGND VPWR VPWR _20302_/A sky130_fd_sc_hd__or3_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21281_ _23685_/Q _20343_/X _23701_/Q _21217_/X VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__o22a_4
X_23020_ _23020_/A _23008_/Y _23013_/X _23020_/D VGND VGND VPWR VPWR _23020_/X sky130_fd_sc_hd__or4_4
X_20232_ _20232_/A VGND VGND VPWR VPWR _20232_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22641__A _22641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20163_ _20150_/Y VGND VGND VPWR VPWR _20163_/X sky130_fd_sc_hd__buf_2
XFILLER_89_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22203__A1 _25531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20094_ _20092_/Y _20093_/X _19734_/X _20093_/X VGND VGND VPWR VPWR _20094_/X sky130_fd_sc_hd__a2bb2o_4
X_24971_ _24975_/CLK _24971_/D HRESETn VGND VGND VPWR VPWR _13908_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11783__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23922_ _25491_/CLK _23922_/D VGND VGND VPWR VPWR _18944_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15255__A _15293_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19080__B1 _19008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24638__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23853_ _23871_/CLK _23853_/D VGND VGND VPWR VPWR _23853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19294__A2_N _19293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22804_ _22479_/A VGND VGND VPWR VPWR _22804_/X sky130_fd_sc_hd__buf_2
XANTENNA__21704__B _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20996_ _20996_/A _20996_/B _20996_/C VGND VGND VPWR VPWR _20997_/A sky130_fd_sc_hd__or3_4
X_23784_ _24252_/CLK _23784_/D VGND VGND VPWR VPWR _23784_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25523_ _25520_/CLK _25523_/D HRESETn VGND VGND VPWR VPWR _25523_/Q sky130_fd_sc_hd__dfrtp_4
X_22735_ _22446_/A _22731_/X _23106_/A _22734_/Y VGND VGND VPWR VPWR _22735_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25454_ _25454_/CLK _25454_/D HRESETn VGND VGND VPWR VPWR _25454_/Q sky130_fd_sc_hd__dfrtp_4
X_22666_ _15718_/A _22665_/X _22148_/C _24838_/Q _22695_/B VGND VGND VPWR VPWR _22666_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22816__A _23148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24405_ _24952_/CLK _24405_/D HRESETn VGND VGND VPWR VPWR _17080_/A sky130_fd_sc_hd__dfrtp_4
X_21617_ _21611_/X _21617_/B _21616_/X VGND VGND VPWR VPWR _21617_/X sky130_fd_sc_hd__and3_4
X_25385_ _25392_/CLK _12947_/Y HRESETn VGND VGND VPWR VPWR _25385_/Q sky130_fd_sc_hd__dfrtp_4
X_22597_ _20885_/Y _21606_/X _20746_/Y _21123_/X VGND VGND VPWR VPWR _22597_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22535__B _22535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _24842_/Q VGND VGND VPWR VPWR _12350_/Y sky130_fd_sc_hd__inv_2
X_24336_ _24337_/CLK _17435_/X HRESETn VGND VGND VPWR VPWR _17432_/A sky130_fd_sc_hd__dfrtp_4
X_21548_ _21090_/A VGND VGND VPWR VPWR _21719_/B sky130_fd_sc_hd__buf_2
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20336__A _20323_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12281_ _12249_/X _12281_/B _12281_/C _12281_/D VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__or4_4
X_21479_ _21470_/X _21478_/X _17732_/X VGND VGND VPWR VPWR _21487_/B sky130_fd_sc_hd__o21a_4
X_24267_ _24715_/CLK _24267_/D HRESETn VGND VGND VPWR VPWR _24267_/Q sky130_fd_sc_hd__dfrtp_4
X_14020_ _13998_/X VGND VGND VPWR VPWR _14020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17236__A1_N _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23218_ _23218_/A _23183_/B VGND VGND VPWR VPWR _23221_/B sky130_fd_sc_hd__or2_4
X_24198_ _24196_/CLK _18392_/X HRESETn VGND VGND VPWR VPWR _24198_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23149_ _24577_/Q _22897_/X _23148_/X VGND VGND VPWR VPWR _23149_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15971_ _12209_/Y _15968_/X _15970_/X _15968_/X VGND VGND VPWR VPWR _24771_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17364__B _17364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17710_ _13781_/A _11718_/B _17455_/X _21178_/A VGND VGND VPWR VPWR _17710_/X sky130_fd_sc_hd__or4_4
X_14922_ _14922_/A VGND VGND VPWR VPWR _14922_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18690_ _18637_/Y _18626_/Y _18614_/Y _18690_/D VGND VGND VPWR VPWR _18690_/X sky130_fd_sc_hd__or4_4
XANTENNA__19071__B1 _19048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17641_ _17641_/A _17639_/X _17640_/X VGND VGND VPWR VPWR _24317_/D sky130_fd_sc_hd__and3_4
XANTENNA__23382__A _21025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14853_ _14834_/X _14851_/Y _25056_/Q _14852_/X VGND VGND VPWR VPWR _14853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _16464_/A _16464_/B _13804_/C _13804_/D VGND VGND VPWR VPWR _13805_/A sky130_fd_sc_hd__and4_4
X_17572_ _17572_/A VGND VGND VPWR VPWR _17573_/A sky130_fd_sc_hd__inv_2
X_14784_ _14773_/Y _14781_/X _25065_/Q _14783_/X VGND VGND VPWR VPWR _14784_/X sky130_fd_sc_hd__o22a_4
X_11996_ _11992_/X VGND VGND VPWR VPWR _11996_/Y sky130_fd_sc_hd__inv_2
X_19311_ _23793_/Q VGND VGND VPWR VPWR _19311_/Y sky130_fd_sc_hd__inv_2
X_16523_ _16522_/Y _16520_/X _16349_/X _16520_/X VGND VGND VPWR VPWR _24562_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13735_ _13693_/X _13734_/Y _13730_/X _13722_/X _11665_/A VGND VGND VPWR VPWR _25290_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19242_ _19240_/Y _19236_/X _19151_/X _19241_/X VGND VGND VPWR VPWR _19242_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21720__A3 _21550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16454_ _24585_/Q VGND VGND VPWR VPWR _16454_/Y sky130_fd_sc_hd__inv_2
X_13666_ _13666_/A _13666_/B VGND VGND VPWR VPWR _13667_/B sky130_fd_sc_hd__or2_4
XFILLER_188_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22726__A _22726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15405_ _15082_/Y _15408_/B _15348_/X VGND VGND VPWR VPWR _15405_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21630__A _21630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12617_ _25427_/Q VGND VGND VPWR VPWR _12679_/A sky130_fd_sc_hd__inv_2
X_19173_ _18062_/B VGND VGND VPWR VPWR _19173_/Y sky130_fd_sc_hd__inv_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ HWDATA[31] VGND VGND VPWR VPWR _16385_/X sky130_fd_sc_hd__buf_2
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13597_ _13597_/A _13573_/X _13587_/X _13596_/X VGND VGND VPWR VPWR _13597_/X sky130_fd_sc_hd__or4_4
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18124_ _17954_/A _18116_/X _18123_/X VGND VGND VPWR VPWR _18124_/X sky130_fd_sc_hd__and3_4
X_15336_ _15336_/A VGND VGND VPWR VPWR _15336_/Y sky130_fd_sc_hd__inv_2
X_12548_ _24884_/Q VGND VGND VPWR VPWR _12548_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18055_ _18231_/A _18055_/B VGND VGND VPWR VPWR _18055_/X sky130_fd_sc_hd__or2_4
X_15267_ _15266_/X VGND VGND VPWR VPWR _25023_/D sky130_fd_sc_hd__inv_2
X_12479_ _12263_/Y _12479_/B VGND VGND VPWR VPWR _12502_/A sky130_fd_sc_hd__or2_4
X_17006_ _16048_/Y _17041_/A _16048_/Y _17041_/A VGND VGND VPWR VPWR _17006_/X sky130_fd_sc_hd__a2bb2o_4
X_14218_ _14218_/A VGND VGND VPWR VPWR _14218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22433__A1 _25380_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15198_ _15080_/B _15181_/B _14910_/Y VGND VGND VPWR VPWR _15198_/X sky130_fd_sc_hd__o21a_4
XFILLER_141_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12159__A1_N _12113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_25_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _24302_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_4_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14149_ _14149_/A VGND VGND VPWR VPWR _14149_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_88_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _24803_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21077__A _21058_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18957_ _18956_/Y _18952_/X _17452_/X _18952_/A VGND VGND VPWR VPWR _18957_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22197__B1 _22185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ _17907_/X VGND VGND VPWR VPWR _17908_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19062__B1 _19012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18888_ _23961_/Q _18888_/B VGND VGND VPWR VPWR _18891_/B sky130_fd_sc_hd__or2_4
XFILLER_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24731__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17839_ _17839_/A VGND VGND VPWR VPWR _24279_/D sky130_fd_sc_hd__inv_2
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _13666_/B VGND VGND VPWR VPWR _20850_/Y sky130_fd_sc_hd__inv_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19509_ _22343_/B _19508_/X _11939_/X _19508_/X VGND VGND VPWR VPWR _23724_/D sky130_fd_sc_hd__a2bb2o_4
X_20781_ _24034_/Q _20776_/X _20780_/Y VGND VGND VPWR VPWR _20781_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__17376__B1 _17280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14419__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22520_ _20735_/Y _21123_/X _20874_/Y _22808_/A VGND VGND VPWR VPWR _22520_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15926__A1 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21540__A _21714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22451_ _22450_/X VGND VGND VPWR VPWR _22451_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21402_ _21398_/X _21402_/B VGND VGND VPWR VPWR _21402_/X sky130_fd_sc_hd__or2_4
X_22382_ _22394_/A _22382_/B VGND VGND VPWR VPWR _22383_/C sky130_fd_sc_hd__or2_4
X_25170_ _25168_/CLK _25170_/D HRESETn VGND VGND VPWR VPWR _12169_/D sky130_fd_sc_hd__dfrtp_4
X_21333_ _21332_/X VGND VGND VPWR VPWR _21591_/A sky130_fd_sc_hd__buf_2
X_24121_ _24121_/CLK MSI_S3 HRESETn VGND VGND VPWR VPWR _24121_/Q sky130_fd_sc_hd__dfrtp_4
X_21264_ _21267_/A _19942_/Y VGND VGND VPWR VPWR _21265_/C sky130_fd_sc_hd__or2_4
X_24052_ _24488_/CLK _20858_/Y HRESETn VGND VGND VPWR VPWR _13666_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_144_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20435__B1 _20249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20215_ _20211_/Y _20214_/X _16866_/X _20214_/X VGND VGND VPWR VPWR _20215_/X sky130_fd_sc_hd__a2bb2o_4
X_23003_ _23003_/A _23140_/B VGND VGND VPWR VPWR _23003_/X sky130_fd_sc_hd__and2_4
XANTENNA__22975__A2 _22531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21195_ _21211_/A _21195_/B VGND VGND VPWR VPWR _21195_/X sky130_fd_sc_hd__or2_4
XFILLER_104_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20146_ _20146_/A VGND VGND VPWR VPWR _20146_/X sky130_fd_sc_hd__buf_2
XANTENNA__24819__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20077_ _21271_/B _20072_/X _19856_/X _20059_/Y VGND VGND VPWR VPWR _20077_/X sky130_fd_sc_hd__a2bb2o_4
X_24954_ _24240_/CLK _24954_/D HRESETn VGND VGND VPWR VPWR _14684_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23905_ _24214_/CLK _23905_/D VGND VGND VPWR VPWR _23905_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21715__A _21715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24885_ _24883_/CLK _15735_/X HRESETn VGND VGND VPWR VPWR _24885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ HWDATA[5] VGND VGND VPWR VPWR _11851_/A sky130_fd_sc_hd__buf_2
X_23836_ _23836_/CLK _19192_/X VGND VGND VPWR VPWR _23836_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11779_/Y _11777_/X _11780_/X _11777_/X VGND VGND VPWR VPWR _25548_/D sky130_fd_sc_hd__a2bb2o_4
X_23767_ _23768_/CLK _19384_/X VGND VGND VPWR VPWR _18142_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21163__A1 _14250_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ _12142_/X _12168_/X VGND VGND VPWR VPWR _20979_/X sky130_fd_sc_hd__and2_4
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _13520_/A VGND VGND VPWR VPWR _13520_/Y sky130_fd_sc_hd__inv_2
X_25506_ _25181_/CLK _11977_/X HRESETn VGND VGND VPWR VPWR _25506_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13233__A _13153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22718_ _24534_/Q _22424_/B _21741_/A _22717_/X VGND VGND VPWR VPWR _22718_/X sky130_fd_sc_hd__a211o_4
XFILLER_213_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23698_ _23408_/CLK _23698_/D VGND VGND VPWR VPWR _23698_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_202_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21450__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13451_ _13451_/A _13449_/X _13451_/C VGND VGND VPWR VPWR _13455_/B sky130_fd_sc_hd__and3_4
X_25437_ _25419_/CLK _25437_/D HRESETn VGND VGND VPWR VPWR _12521_/A sky130_fd_sc_hd__dfrtp_4
X_22649_ _22649_/A _23053_/A VGND VGND VPWR VPWR _22649_/X sky130_fd_sc_hd__or2_4
XFILLER_167_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12402_ _12282_/X VGND VGND VPWR VPWR _12403_/A sky130_fd_sc_hd__inv_2
X_16170_ _16169_/Y _16167_/X _15483_/X _16167_/X VGND VGND VPWR VPWR _24689_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22663__A1 _15718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13382_ _13222_/X _23455_/Q VGND VGND VPWR VPWR _13382_/X sky130_fd_sc_hd__or2_4
X_25368_ _25368_/CLK _13028_/Y HRESETn VGND VGND VPWR VPWR _12994_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17359__B _17364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18867__B1 _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22663__B2 _16003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _15121_/A VGND VGND VPWR VPWR _15121_/Y sky130_fd_sc_hd__inv_2
X_12333_ _24832_/Q VGND VGND VPWR VPWR _12333_/Y sky130_fd_sc_hd__inv_2
X_24319_ _24327_/CLK _17630_/X HRESETn VGND VGND VPWR VPWR _24319_/Q sky130_fd_sc_hd__dfrtp_4
X_25299_ _24406_/CLK _13713_/X HRESETn VGND VGND VPWR VPWR _11705_/A sky130_fd_sc_hd__dfrtp_4
X_15052_ _14927_/A _15051_/Y _14927_/A _15051_/Y VGND VGND VPWR VPWR _15052_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22415__A1 _25532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23377__A _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12264_ _23228_/A VGND VGND VPWR VPWR _12264_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_241_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24145_/CLK sky130_fd_sc_hd__clkbuf_1
X_14003_ _14003_/A VGND VGND VPWR VPWR _14003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20426__B1 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17375__A _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12195_ _12187_/X _12189_/X _12192_/X _12195_/D VGND VGND VPWR VPWR _12236_/A sky130_fd_sc_hd__or4_4
X_19860_ _19859_/X _13771_/X _19278_/X VGND VGND VPWR VPWR _19861_/A sky130_fd_sc_hd__or3_4
XFILLER_150_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18811_ _18630_/Y _18810_/X _18714_/X VGND VGND VPWR VPWR _18811_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16812__A2_N _16806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19791_ _19786_/Y _19789_/X _19790_/X _19789_/X VGND VGND VPWR VPWR _23628_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22718__A2 _22424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15954_ _12203_/Y _15947_/X _15952_/X _15953_/X VGND VGND VPWR VPWR _15954_/X sky130_fd_sc_hd__a2bb2o_4
X_18742_ _18742_/A VGND VGND VPWR VPWR _18742_/Y sky130_fd_sc_hd__inv_2
X_14905_ _14905_/A _14898_/X _14901_/X _14904_/X VGND VGND VPWR VPWR _14905_/X sky130_fd_sc_hd__or4_4
XFILLER_37_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18673_ _18673_/A _18673_/B _18673_/C _18672_/X VGND VGND VPWR VPWR _18673_/X sky130_fd_sc_hd__or4_4
X_15885_ _15858_/X _15865_/X _15738_/X _23054_/A _15872_/X VGND VGND VPWR VPWR _24813_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15605__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ _14806_/A _14812_/X _14806_/Y _14815_/B VGND VGND VPWR VPWR _14836_/X sky130_fd_sc_hd__o22a_4
X_17624_ _17573_/A _17627_/B _17600_/X VGND VGND VPWR VPWR _17624_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19124__A2_N _19121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17555_ _17548_/X _17555_/B _17552_/X _17554_/X VGND VGND VPWR VPWR _17555_/X sky130_fd_sc_hd__or4_4
X_14767_ _14766_/X VGND VGND VPWR VPWR _21629_/A sky130_fd_sc_hd__buf_2
XANTENNA__21154__A1 _12132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11979_ _11979_/A _11979_/B _11979_/C _11712_/B VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__or4_4
X_16506_ _16506_/A VGND VGND VPWR VPWR _16506_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13718_ _13707_/B _13716_/X _13717_/Y _13712_/X _11666_/A VGND VGND VPWR VPWR _25297_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ _17485_/Y _17459_/A VGND VGND VPWR VPWR _17486_/X sky130_fd_sc_hd__or2_4
X_14698_ _21914_/A VGND VGND VPWR VPWR _14761_/A sky130_fd_sc_hd__buf_2
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16437_ _15095_/Y _16435_/X _16349_/X _16435_/X VGND VGND VPWR VPWR _24595_/D sky130_fd_sc_hd__a2bb2o_4
X_19225_ _19225_/A VGND VGND VPWR VPWR _19225_/X sky130_fd_sc_hd__buf_2
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13649_ _13535_/Y VGND VGND VPWR VPWR _13649_/X sky130_fd_sc_hd__buf_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16454__A _24585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19156_ _23848_/Q VGND VGND VPWR VPWR _19156_/Y sky130_fd_sc_hd__inv_2
X_16368_ _14412_/A VGND VGND VPWR VPWR _16368_/X sky130_fd_sc_hd__buf_2
XFILLER_185_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18107_ _18107_/A _18107_/B _18107_/C VGND VGND VPWR VPWR _18107_/X sky130_fd_sc_hd__and3_4
XFILLER_145_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_51_0_HCLK clkbuf_6_50_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15319_ _15164_/Y _15337_/A _15318_/X VGND VGND VPWR VPWR _15319_/X sky130_fd_sc_hd__or3_4
X_19087_ _13346_/B VGND VGND VPWR VPWR _19087_/Y sky130_fd_sc_hd__inv_2
X_16299_ _16296_/Y _16291_/X _15948_/X _16298_/X VGND VGND VPWR VPWR _24646_/D sky130_fd_sc_hd__a2bb2o_4
X_18038_ _18006_/A VGND VGND VPWR VPWR _18039_/A sky130_fd_sc_hd__buf_2
XFILLER_172_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20000_ _20000_/A VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__buf_2
XANTENNA__20968__B2 _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24912__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19989_ _19988_/Y VGND VGND VPWR VPWR _19989_/X sky130_fd_sc_hd__buf_2
XANTENNA__14647__A1 _13547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19035__B1 _19008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21535__A _21535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21951_ _21679_/A _21940_/X _21950_/X VGND VGND VPWR VPWR _21951_/X sky130_fd_sc_hd__or3_4
XFILLER_223_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16629__A _24521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20902_ _20907_/B VGND VGND VPWR VPWR _20911_/B sky130_fd_sc_hd__inv_2
XFILLER_27_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15533__A _15544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24670_ _24552_/CLK _16230_/X HRESETn VGND VGND VPWR VPWR _16229_/A sky130_fd_sc_hd__dfrtp_4
X_21882_ _21882_/A VGND VGND VPWR VPWR _22954_/C sky130_fd_sc_hd__buf_2
XFILLER_242_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23445_/CLK _19813_/X VGND VGND VPWR VPWR _19812_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20854_/A VGND VGND VPWR VPWR _20833_/X sky130_fd_sc_hd__buf_2
XFILLER_242_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22342__B1 _22329_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23552_ _23553_/CLK _20004_/X VGND VGND VPWR VPWR _20002_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20764_ _13142_/C _20758_/X _20763_/Y VGND VGND VPWR VPWR _20764_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12830__B1 _25401_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _21445_/X VGND VGND VPWR VPWR _22503_/X sky130_fd_sc_hd__buf_2
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _20716_/A VGND VGND VPWR VPWR _20695_/X sky130_fd_sc_hd__buf_2
X_23483_ _23516_/CLK _23483_/D VGND VGND VPWR VPWR _20195_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25222_ _25223_/CLK _25222_/D HRESETn VGND VGND VPWR VPWR _14124_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22434_ _23299_/A _22427_/Y _22430_/X _22431_/X _22433_/X VGND VGND VPWR VPWR _22435_/D
+ sky130_fd_sc_hd__o32a_4
XANTENNA__18849__B1 _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25203__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25153_ _24334_/CLK _25153_/D HRESETn VGND VGND VPWR VPWR _25153_/Q sky130_fd_sc_hd__dfrtp_4
X_22365_ _21476_/A _22365_/B VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__or2_4
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24104_ _23631_/CLK _24104_/D HRESETn VGND VGND VPWR VPWR _12000_/B sky130_fd_sc_hd__dfrtp_4
X_21316_ _22577_/B VGND VGND VPWR VPWR _21316_/X sky130_fd_sc_hd__buf_2
X_22296_ _21606_/A VGND VGND VPWR VPWR _22296_/X sky130_fd_sc_hd__buf_2
X_25084_ _25062_/CLK _14644_/X HRESETn VGND VGND VPWR VPWR _14626_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22948__A2 _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21247_ _21273_/A _21247_/B VGND VGND VPWR VPWR _21250_/B sky130_fd_sc_hd__or2_4
X_24035_ _24500_/CLK _20787_/X HRESETn VGND VGND VPWR VPWR _20790_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_151_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20959__B2 _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24653__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21178_ _21178_/A VGND VGND VPWR VPWR _21967_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_71_0_HCLK clkbuf_8_70_0_HCLK/A VGND VGND VPWR VPWR _24792_/CLK sky130_fd_sc_hd__clkbuf_1
X_20129_ _20129_/A VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13228__A _13228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12649__B1 _12657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12951_ _12828_/X _12950_/X VGND VGND VPWR VPWR _12952_/D sky130_fd_sc_hd__or2_4
X_24937_ _24937_/CLK _15539_/X HRESETn VGND VGND VPWR VPWR _21135_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15850__A3 _15782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15546__A1_N _12107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16539__A _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22581__B1 _21844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _11902_/A VGND VGND VPWR VPWR _11902_/Y sky130_fd_sc_hd__inv_2
X_15670_ _21031_/A _13821_/B VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__or2_4
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12882_ _12906_/A _12880_/X _12881_/X VGND VGND VPWR VPWR _25402_/D sky130_fd_sc_hd__and3_4
X_24868_ _24867_/CLK _15769_/X HRESETn VGND VGND VPWR VPWR _12545_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16260__B1 _16157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _13593_/A _14608_/X _13779_/X _14569_/B VGND VGND VPWR VPWR _25088_/D sky130_fd_sc_hd__o22a_4
XPHY_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _25534_/Q VGND VGND VPWR VPWR _11833_/Y sky130_fd_sc_hd__inv_2
X_23819_ _23459_/CLK _23819_/D VGND VGND VPWR VPWR _13220_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _24799_/CLK _15907_/X HRESETn VGND VGND VPWR VPWR _22490_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17340_/A _17340_/B VGND VGND VPWR VPWR _17342_/B sky130_fd_sc_hd__or2_4
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _14059_/B _14060_/B VGND VGND VPWR VPWR _14552_/X sky130_fd_sc_hd__or3_4
XFILLER_187_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11762_/Y _11760_/X _11763_/X _11760_/X VGND VGND VPWR VPWR _11764_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13502_/Y _13498_/X _13481_/X _13486_/A VGND VGND VPWR VPWR _13503_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17271_/A VGND VGND VPWR VPWR _17271_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _25126_/Q VGND VGND VPWR VPWR _14483_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _24239_/Q VGND VGND VPWR VPWR _11695_/Y sky130_fd_sc_hd__inv_2
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _23898_/Q VGND VGND VPWR VPWR _19010_/Y sky130_fd_sc_hd__inv_2
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _16227_/A VGND VGND VPWR VPWR _16222_/X sky130_fd_sc_hd__buf_2
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13217_/X _13432_/X _13434_/C VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__and3_4
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16153_ HWDATA[9] VGND VGND VPWR VPWR _16153_/X sky130_fd_sc_hd__buf_2
X_13365_ _13257_/X _13365_/B VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__or2_4
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15104_ _25000_/Q VGND VGND VPWR VPWR _15305_/A sky130_fd_sc_hd__inv_2
XFILLER_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12316_ _25350_/Q _12314_/Y _13026_/A _24851_/Q VGND VGND VPWR VPWR _12316_/X sky130_fd_sc_hd__a2bb2o_4
X_16084_ _24721_/Q VGND VGND VPWR VPWR _16084_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15669__A3 _15656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13296_ _13320_/A VGND VGND VPWR VPWR _13369_/A sky130_fd_sc_hd__buf_2
XFILLER_181_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15035_ _15232_/A _24468_/Q _14912_/X _15034_/Y VGND VGND VPWR VPWR _15035_/X sky130_fd_sc_hd__a2bb2o_4
X_19912_ _23585_/Q VGND VGND VPWR VPWR _21955_/B sky130_fd_sc_hd__inv_2
XFILLER_142_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _12247_/A VGND VGND VPWR VPWR _12247_/X sky130_fd_sc_hd__buf_2
XANTENNA__16079__B1 _15483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _19843_/A VGND VGND VPWR VPWR _19843_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12178_ _12132_/Y _12177_/Y SCLK_S3 _12177_/A VGND VGND VPWR VPWR _12178_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19774_ _19771_/Y _19766_/X _19772_/X _19773_/X VGND VGND VPWR VPWR _23634_/D sky130_fd_sc_hd__a2bb2o_4
X_16986_ _24745_/Q _24402_/Q _16023_/Y _17088_/A VGND VGND VPWR VPWR _16989_/C sky130_fd_sc_hd__o22a_4
XFILLER_84_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18725_ _18727_/B VGND VGND VPWR VPWR _18725_/Y sky130_fd_sc_hd__inv_2
X_15937_ _15678_/X _15796_/X _15933_/X _24785_/Q _15936_/X VGND VGND VPWR VPWR _15937_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22572__B1 _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15868_ _23053_/A VGND VGND VPWR VPWR _21069_/B sky130_fd_sc_hd__buf_2
X_18656_ _16588_/Y _18768_/A _16578_/A _18756_/A VGND VGND VPWR VPWR _18659_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14819_ _14837_/A VGND VGND VPWR VPWR _14819_/X sky130_fd_sc_hd__buf_2
X_17607_ _17525_/Y _17604_/X VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__or2_4
X_15799_ _21043_/A VGND VGND VPWR VPWR _15800_/A sky130_fd_sc_hd__buf_2
X_18587_ _18567_/X VGND VGND VPWR VPWR _18588_/B sky130_fd_sc_hd__inv_2
X_17538_ _17538_/A VGND VGND VPWR VPWR _17588_/A sky130_fd_sc_hd__inv_2
XFILLER_189_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19078__A2_N _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17469_ _17478_/B VGND VGND VPWR VPWR _18333_/C sky130_fd_sc_hd__buf_2
XANTENNA__15800__B _15934_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16184__A _13599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19208_ _19207_/Y _19203_/X _19139_/X _19196_/A VGND VGND VPWR VPWR _23829_/D sky130_fd_sc_hd__a2bb2o_4
X_20480_ _14395_/Y _14504_/X _24095_/Q VGND VGND VPWR VPWR _20480_/X sky130_fd_sc_hd__a21o_4
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19139_ _19139_/A VGND VGND VPWR VPWR _19139_/X sky130_fd_sc_hd__buf_2
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22150_ _22150_/A _22149_/X VGND VGND VPWR VPWR _22150_/X sky130_fd_sc_hd__and2_4
XFILLER_145_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21101_ _22533_/A VGND VGND VPWR VPWR _21101_/X sky130_fd_sc_hd__buf_2
XFILLER_172_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22081_ _21259_/A VGND VGND VPWR VPWR _22394_/A sky130_fd_sc_hd__buf_2
X_21032_ _21031_/X _21577_/A _13822_/A _21045_/A VGND VGND VPWR VPWR _21032_/X sky130_fd_sc_hd__or4_4
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15247__B _15294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15817__B1 _11783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_58_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__24064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15832__A3 _15759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17462__B _17461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _22777_/X _22982_/X _22872_/X _12317_/A _22779_/X VGND VGND VPWR VPWR _22983_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24722_ _24726_/CLK _16083_/X HRESETn VGND VGND VPWR VPWR _24722_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21934_ _21949_/A _21931_/X _21933_/X VGND VGND VPWR VPWR _21934_/X sky130_fd_sc_hd__and3_4
XFILLER_227_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24653_ _24169_/CLK _24653_/D HRESETn VGND VGND VPWR VPWR _21340_/A sky130_fd_sc_hd__dfrtp_4
X_21865_ _12009_/Y _12107_/X _12045_/Y _12080_/X VGND VGND VPWR VPWR _21865_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _25068_/CLK _19863_/X VGND VGND VPWR VPWR _23604_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_24_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20815_/X VGND VGND VPWR VPWR _20816_/Y sky130_fd_sc_hd__inv_2
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24584_ _24657_/CLK _24584_/D HRESETn VGND VGND VPWR VPWR _24584_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12803__B1 _12952_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21712__B _23016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21796_ _19610_/A _21971_/B _23704_/Q _21656_/X VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__o22a_4
XFILLER_242_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18293__B _17712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20609__A _20609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _23590_/CLK _20052_/X VGND VGND VPWR VPWR _20050_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15710__B _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20747_ _20746_/Y _20740_/Y _13140_/X VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__o21a_4
XFILLER_196_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16094__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23466_ _23466_/CLK _23466_/D VGND VGND VPWR VPWR _23466_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15899__A3 _16241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20678_ _20677_/X VGND VGND VPWR VPWR _20678_/Y sky130_fd_sc_hd__inv_2
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25205_ _23998_/CLK _25205_/D HRESETn VGND VGND VPWR VPWR _25205_/Q sky130_fd_sc_hd__dfstp_4
X_22417_ _21511_/X _18278_/X _22410_/X _22415_/X _22416_/X VGND VGND VPWR VPWR _22435_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23291__A1 _21881_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23397_ _24206_/CLK _20417_/X VGND VGND VPWR VPWR _23397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13150_ _13150_/A VGND VGND VPWR VPWR _13150_/Y sky130_fd_sc_hd__inv_2
X_25136_ _25148_/CLK _25136_/D HRESETn VGND VGND VPWR VPWR _25136_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__24834__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22348_ _21945_/A _22348_/B _22348_/C VGND VGND VPWR VPWR _22348_/X sky130_fd_sc_hd__and3_4
XFILLER_136_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12101_ _25483_/Q VGND VGND VPWR VPWR _12101_/Y sky130_fd_sc_hd__inv_2
X_13081_ _13006_/B _13080_/X VGND VGND VPWR VPWR _13084_/B sky130_fd_sc_hd__or2_4
X_25067_ _25066_/CLK _14763_/X HRESETn VGND VGND VPWR VPWR _14687_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19247__B1 _19246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22279_ _21278_/X _22259_/X _22274_/X _22277_/Y _22278_/X VGND VGND VPWR VPWR _22279_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_105_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12334__A2 _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12032_ _12032_/A VGND VGND VPWR VPWR _12032_/Y sky130_fd_sc_hd__inv_2
X_24018_ _24485_/CLK _20711_/Y HRESETn VGND VGND VPWR VPWR _24018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_239_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17653__A _17578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16840_ _16838_/Y _16834_/X _15754_/X _16839_/X VGND VGND VPWR VPWR _16840_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15284__A1 _15258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16481__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23346__A2 _22673_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16771_ _16770_/Y _16768_/X _15752_/X _16768_/X VGND VGND VPWR VPWR _24466_/D sky130_fd_sc_hd__a2bb2o_4
X_13983_ _25247_/Q VGND VGND VPWR VPWR _13984_/A sky130_fd_sc_hd__inv_2
XANTENNA__12797__A _21537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15722_ _15713_/X VGND VGND VPWR VPWR _15722_/X sky130_fd_sc_hd__buf_2
X_18510_ _18510_/A _18510_/B VGND VGND VPWR VPWR _18510_/X sky130_fd_sc_hd__or2_4
XANTENNA__15173__A _15172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ _12933_/X VGND VGND VPWR VPWR _12934_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19490_ _22038_/B _19484_/X _11948_/X _19489_/X VGND VGND VPWR VPWR _19490_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15653_ _15653_/A _11740_/C _11740_/D _14442_/A VGND VGND VPWR VPWR _15657_/A sky130_fd_sc_hd__or4_4
X_18441_ _16231_/Y _24180_/Q _24673_/Q _18534_/A VGND VGND VPWR VPWR _18443_/C sky130_fd_sc_hd__a2bb2o_4
X_12865_ _12638_/B _12872_/A VGND VGND VPWR VPWR _12865_/X sky130_fd_sc_hd__or2_4
XFILLER_46_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14577_/B _14595_/X _14603_/Y _14599_/X _25096_/Q VGND VGND VPWR VPWR _14604_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_221_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11816_/A VGND VGND VPWR VPWR _11816_/Y sky130_fd_sc_hd__inv_2
X_18372_ _18372_/A _18358_/X VGND VGND VPWR VPWR _18372_/X sky130_fd_sc_hd__or2_4
XPHY_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/A VGND VGND VPWR VPWR _15584_/X sky130_fd_sc_hd__buf_2
XFILLER_187_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _25375_/Q VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__inv_2
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17315_/X _17321_/X _17323_/C VGND VGND VPWR VPWR _24367_/D sky130_fd_sc_hd__and3_4
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _25110_/Q _14519_/X _21560_/A _14514_/X VGND VGND VPWR VPWR _14535_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11747_/A VGND VGND VPWR VPWR _22694_/B sky130_fd_sc_hd__buf_2
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17254_ _17253_/Y _17389_/A _17214_/Y VGND VGND VPWR VPWR _17255_/D sky130_fd_sc_hd__or3_4
XFILLER_186_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14465_/Y _14463_/X _14423_/X _14463_/X VGND VGND VPWR VPWR _25133_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _11678_/A VGND VGND VPWR VPWR _13736_/A sky130_fd_sc_hd__inv_2
XFILLER_174_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16205_ _23250_/A VGND VGND VPWR VPWR _16205_/Y sky130_fd_sc_hd__inv_2
X_13417_ _13417_/A _23934_/Q VGND VGND VPWR VPWR _13417_/X sky130_fd_sc_hd__or2_4
X_17185_ _16348_/A _17359_/C _16304_/Y _17245_/A VGND VGND VPWR VPWR _17185_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23282__A1 _16102_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14397_ _20438_/A VGND VGND VPWR VPWR _20470_/A sky130_fd_sc_hd__inv_2
XANTENNA__16732__A _16731_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24100__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16136_ _16162_/A VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__buf_2
XANTENNA__24575__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13348_ _13412_/A _13346_/X _13348_/C VGND VGND VPWR VPWR _13352_/B sky130_fd_sc_hd__and3_4
XFILLER_155_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11781__B1 _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11876__A _13481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _16065_/Y _16061_/X _16066_/X _16061_/X VGND VGND VPWR VPWR _24728_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ _13317_/A _18965_/A VGND VGND VPWR VPWR _13280_/C sky130_fd_sc_hd__or2_4
XFILLER_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21069__B _21069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15018_ _14924_/A _15017_/A _15268_/A _15017_/Y VGND VGND VPWR VPWR _15021_/C sky130_fd_sc_hd__o22a_4
XFILLER_142_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12325__A2 _24844_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19826_ _23616_/Q VGND VGND VPWR VPWR _19826_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17563__A _17562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__A3 _15734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21085__A _21085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19757_ _19755_/Y _19756_/X _19734_/X _19756_/X VGND VGND VPWR VPWR _19757_/X sky130_fd_sc_hd__a2bb2o_4
X_16969_ _24384_/Q VGND VGND VPWR VPWR _16969_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18708_ _18606_/X _18708_/B VGND VGND VPWR VPWR _18709_/C sky130_fd_sc_hd__nand2_4
XFILLER_65_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19688_ _13393_/B VGND VGND VPWR VPWR _19688_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18639_ _24529_/Q _24140_/Q _16608_/Y _18805_/A VGND VGND VPWR VPWR _18639_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21650_ _21646_/X _21649_/X _14758_/X VGND VGND VPWR VPWR _21650_/X sky130_fd_sc_hd__o21a_4
XFILLER_212_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20601_ _18888_/B VGND VGND VPWR VPWR _20601_/Y sky130_fd_sc_hd__inv_2
X_21581_ _13520_/Y _21579_/X _12049_/Y _21580_/X VGND VGND VPWR VPWR _21581_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14427__A _14427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23320_ _21547_/X _23319_/X _23159_/X _24856_/Q _22851_/X VGND VGND VPWR VPWR _23320_/X
+ sky130_fd_sc_hd__a32o_4
X_20532_ _24088_/Q _24093_/Q _24089_/Q VGND VGND VPWR VPWR _20532_/X sky130_fd_sc_hd__or3_4
XFILLER_192_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22644__A _22644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20463_ _20463_/A _20445_/A _20463_/C VGND VGND VPWR VPWR _20463_/X sky130_fd_sc_hd__and3_4
X_23251_ _16478_/A _23184_/X _23148_/X VGND VGND VPWR VPWR _23251_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12357__A2_N _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22202_ _21877_/B _22202_/B _22202_/C VGND VGND VPWR VPWR _22202_/X sky130_fd_sc_hd__and3_4
Xclkbuf_5_21_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20394_ _21952_/B _20391_/X _19636_/A _20391_/X VGND VGND VPWR VPWR _23408_/D sky130_fd_sc_hd__a2bb2o_4
X_23182_ _23249_/A _23181_/X VGND VGND VPWR VPWR _23182_/Y sky130_fd_sc_hd__nor2_4
XFILLER_192_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22481__C1 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _22132_/X VGND VGND VPWR VPWR _22133_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15258__A _15258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19229__B1 _19184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22064_ _19605_/Y _19597_/X VGND VGND VPWR VPWR _22064_/X sky130_fd_sc_hd__and2_4
XFILLER_87_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21587__A1 _21565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21015_ _21014_/X VGND VGND VPWR VPWR _21015_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15805__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_145_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _25309_/CLK sky130_fd_sc_hd__clkbuf_1
X_22966_ _22966_/A VGND VGND VPWR VPWR _22966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22819__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15018__B2 _15017_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24705_ _25444_/CLK _24705_/D HRESETn VGND VGND VPWR VPWR _22920_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21917_ _21914_/A _21917_/B VGND VGND VPWR VPWR _21919_/B sky130_fd_sc_hd__or2_4
XFILLER_215_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22897_ _22897_/A VGND VGND VPWR VPWR _22897_/X sky130_fd_sc_hd__buf_2
XFILLER_71_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12650_ _12649_/X VGND VGND VPWR VPWR _12650_/Y sky130_fd_sc_hd__inv_2
X_24636_ _24629_/CLK _24636_/D HRESETn VGND VGND VPWR VPWR _24636_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21848_ _21847_/Y _21161_/X _17436_/Y _17424_/X VGND VGND VPWR VPWR _21848_/X sky130_fd_sc_hd__o22a_4
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _25429_/Q VGND VGND VPWR VPWR _12660_/A sky130_fd_sc_hd__inv_2
X_24567_ _24601_/CLK _24567_/D HRESETn VGND VGND VPWR VPWR _16510_/A sky130_fd_sc_hd__dfrtp_4
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21779_ _22388_/A _20181_/Y VGND VGND VPWR VPWR _21781_/B sky130_fd_sc_hd__or2_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _14320_/A VGND VGND VPWR VPWR _14320_/X sky130_fd_sc_hd__buf_2
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23518_ _23918_/CLK _20096_/X VGND VGND VPWR VPWR _20095_/A sky130_fd_sc_hd__dfxtp_4
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24498_ _24532_/CLK _16695_/X HRESETn VGND VGND VPWR VPWR _24498_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16783__A1_N _15022_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14250_/Y _14245_/X _13819_/X _14233_/A VGND VGND VPWR VPWR _14251_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _23529_/CLK _23449_/D VGND VGND VPWR VPWR _23449_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16552__A _16552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _13187_/X _13194_/X _13201_/X _11979_/A _11979_/C VGND VGND VPWR VPWR _13202_/X
+ sky130_fd_sc_hd__o32a_4
X_14182_ _14174_/B _14181_/X VGND VGND VPWR VPWR _14182_/Y sky130_fd_sc_hd__nor2_4
XFILLER_152_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16168__A1_N _16166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13133_ _13132_/X VGND VGND VPWR VPWR _13134_/B sky130_fd_sc_hd__inv_2
X_25119_ _25154_/CLK _25119_/D HRESETn VGND VGND VPWR VPWR _25119_/Q sky130_fd_sc_hd__dfrtp_4
X_18990_ _23904_/Q VGND VGND VPWR VPWR _18990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16798__A1_N _15019_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13064_ _12323_/Y _13069_/B _13040_/X VGND VGND VPWR VPWR _13064_/Y sky130_fd_sc_hd__a21oi_4
X_17941_ _17941_/A _17939_/X _17940_/X VGND VGND VPWR VPWR _17941_/X sky130_fd_sc_hd__and3_4
X_12015_ _12015_/A VGND VGND VPWR VPWR _12015_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17872_ _17861_/A _17872_/B VGND VGND VPWR VPWR _17873_/C sky130_fd_sc_hd__or2_4
XFILLER_239_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19611_ _19610_/X VGND VGND VPWR VPWR _19611_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_41_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16823_ _16822_/Y _16820_/X _15738_/X _16820_/X VGND VGND VPWR VPWR _24442_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19542_ _21692_/B _19541_/X _11961_/X _19541_/X VGND VGND VPWR VPWR _23711_/D sky130_fd_sc_hd__a2bb2o_4
X_13966_ _24980_/Q _13942_/X VGND VGND VPWR VPWR _13967_/B sky130_fd_sc_hd__or2_4
X_16754_ _16754_/A VGND VGND VPWR VPWR _16754_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16206__B1 _15950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22729__A _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12917_ _12857_/Y _12917_/B VGND VGND VPWR VPWR _12918_/C sky130_fd_sc_hd__or2_4
X_15705_ _15696_/A _15696_/B _15704_/X VGND VGND VPWR VPWR _15705_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19943__B2 _19925_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16685_ _16685_/A VGND VGND VPWR VPWR _16685_/X sky130_fd_sc_hd__buf_2
X_19473_ _19460_/Y VGND VGND VPWR VPWR _19473_/X sky130_fd_sc_hd__buf_2
XFILLER_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13897_ _24980_/Q VGND VGND VPWR VPWR _13944_/A sky130_fd_sc_hd__buf_2
X_18424_ _24661_/Q _18423_/A _16256_/Y _18476_/A VGND VGND VPWR VPWR _18424_/X sky130_fd_sc_hd__o22a_4
X_12848_ _12988_/A VGND VGND VPWR VPWR _12906_/A sky130_fd_sc_hd__buf_2
X_15636_ _14427_/A VGND VGND VPWR VPWR _15636_/X sky130_fd_sc_hd__buf_2
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20249__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15567_ _15557_/X _15561_/Y _15562_/X _23336_/A _15569_/A VGND VGND VPWR VPWR _24929_/D
+ sky130_fd_sc_hd__a32o_4
X_18355_ _24206_/Q VGND VGND VPWR VPWR _18355_/Y sky130_fd_sc_hd__inv_2
X_12779_ _25381_/Q _24798_/Q _12777_/X _12778_/Y VGND VGND VPWR VPWR _12779_/X sky130_fd_sc_hd__o22a_4
XFILLER_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _25116_/Q _14516_/X _14524_/A _14517_/Y VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__a211o_4
X_17306_ _17242_/X _17304_/X _17306_/C VGND VGND VPWR VPWR _24371_/D sky130_fd_sc_hd__and3_4
XFILLER_175_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24756__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15498_ _15497_/X VGND VGND VPWR VPWR _15499_/A sky130_fd_sc_hd__inv_2
X_18286_ _17733_/A VGND VGND VPWR VPWR _18286_/Y sky130_fd_sc_hd__inv_2
X_14449_ _14448_/Y _14446_/X _14423_/X _14446_/X VGND VGND VPWR VPWR _25141_/D sky130_fd_sc_hd__a2bb2o_4
X_17237_ _16358_/Y _17177_/A _16367_/Y _17253_/A VGND VGND VPWR VPWR _17238_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17168_ _17137_/B _17163_/X VGND VGND VPWR VPWR _17168_/Y sky130_fd_sc_hd__nand2_4
XFILLER_162_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16119_ _16118_/Y _16116_/X _11780_/X _16116_/X VGND VGND VPWR VPWR _24709_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19773__A _19765_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17099_ _17064_/A VGND VGND VPWR VPWR _17106_/A sky130_fd_sc_hd__buf_2
XANTENNA__23007__B2 _21229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16693__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15930__A1_N _15694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21808__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15806__A _15826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19809_ _23622_/Q VGND VGND VPWR VPWR _19809_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22820_ _24668_/Q _15681_/X VGND VGND VPWR VPWR _22823_/B sky130_fd_sc_hd__or2_4
XFILLER_226_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12230__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_218_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24542_/CLK sky130_fd_sc_hd__clkbuf_1
X_22751_ _22751_/A _22589_/B VGND VGND VPWR VPWR _22754_/B sky130_fd_sc_hd__or2_4
XFILLER_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21702_ _13804_/D _21701_/X _18273_/A _18268_/X VGND VGND VPWR VPWR _21702_/X sky130_fd_sc_hd__o22a_4
XFILLER_212_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25470_ _24196_/CLK _25470_/D HRESETn VGND VGND VPWR VPWR _12184_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19013__A _19020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22682_ _22682_/A _21882_/A VGND VGND VPWR VPWR _22682_/X sky130_fd_sc_hd__and2_4
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24421_ _24613_/CLK _16862_/X HRESETn VGND VGND VPWR VPWR _24421_/Q sky130_fd_sc_hd__dfrtp_4
X_21633_ _21257_/A VGND VGND VPWR VPWR _22388_/A sky130_fd_sc_hd__buf_2
XFILLER_178_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20229__A2_N _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24625_/CLK _17379_/X HRESETn VGND VGND VPWR VPWR _17177_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12785__A2 _22428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21564_ _21731_/A _21564_/B VGND VGND VPWR VPWR _21564_/Y sky130_fd_sc_hd__nor2_4
XFILLER_178_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23303_ _23303_/A _23303_/B VGND VGND VPWR VPWR _23303_/X sky130_fd_sc_hd__and2_4
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20515_ _14395_/A _14504_/X _20513_/X _20477_/C _20514_/X VGND VGND VPWR VPWR _20515_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15184__B1 _15183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24283_ _24283_/CLK _17827_/Y HRESETn VGND VGND VPWR VPWR _16950_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21495_ _21687_/A _21495_/B VGND VGND VPWR VPWR _21498_/B sky130_fd_sc_hd__or2_4
XFILLER_153_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23234_ _24645_/Q _21536_/X VGND VGND VPWR VPWR _23234_/X sky130_fd_sc_hd__or2_4
X_20446_ _13985_/X _20613_/A _20446_/C _20445_/X VGND VGND VPWR VPWR _20446_/X sky130_fd_sc_hd__or4_4
XFILLER_165_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16091__B _15683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23165_ _24643_/Q _23165_/B VGND VGND VPWR VPWR _23165_/X sky130_fd_sc_hd__or2_4
X_20377_ _20364_/Y VGND VGND VPWR VPWR _20377_/X sky130_fd_sc_hd__buf_2
X_22116_ _22115_/Y _21353_/X _14425_/Y _21356_/X VGND VGND VPWR VPWR _22117_/A sky130_fd_sc_hd__o22a_4
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21718__A _21126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23096_ _20944_/B _21306_/A _13145_/B _21607_/X VGND VGND VPWR VPWR _23096_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__18299__A _21210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22047_ _22028_/A _22047_/B VGND VGND VPWR VPWR _22047_/X sky130_fd_sc_hd__or2_4
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16436__B1 _16252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22509__B1 _12793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _13817_/Y _13813_/X _13819_/X _13813_/X VGND VGND VPWR VPWR _25276_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13236__A _13320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23998_ _23998_/CLK _20675_/X HRESETn VGND VGND VPWR VPWR _17407_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13751_ _14775_/B VGND VGND VPWR VPWR _13751_/Y sky130_fd_sc_hd__inv_2
X_22949_ _14936_/A _22947_/X _22542_/A _22948_/X VGND VGND VPWR VPWR _22950_/C sky130_fd_sc_hd__a211o_4
XFILLER_44_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12702_ _12702_/A _12626_/X VGND VGND VPWR VPWR _12702_/X sky130_fd_sc_hd__or2_4
XFILLER_232_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16470_ _16469_/X VGND VGND VPWR VPWR _16470_/X sky130_fd_sc_hd__buf_2
XANTENNA__21172__B _21172_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13682_ _13654_/X VGND VGND VPWR VPWR _13682_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15421_ _15153_/Y _15397_/X _15419_/B _15348_/X VGND VGND VPWR VPWR _15421_/X sky130_fd_sc_hd__a211o_4
XFILLER_203_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12633_ _12633_/A VGND VGND VPWR VPWR _12633_/Y sky130_fd_sc_hd__inv_2
X_24619_ _24625_/CLK _16371_/X HRESETn VGND VGND VPWR VPWR _24619_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20299__A1 _23444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15352_ _15355_/A _15352_/B _15351_/Y VGND VGND VPWR VPWR _25005_/D sky130_fd_sc_hd__and3_4
X_18140_ _15704_/X _18124_/X _18139_/X _24251_/Q _18029_/X VGND VGND VPWR VPWR _18140_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _24878_/Q VGND VGND VPWR VPWR _12564_/Y sky130_fd_sc_hd__inv_2
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22284__A _21450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _14303_/A _14303_/B VGND VGND VPWR VPWR _14304_/A sky130_fd_sc_hd__or2_4
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18071_ _17973_/X _18070_/X _24252_/Q _18031_/X VGND VGND VPWR VPWR _18071_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ _15255_/X _15276_/B _15283_/C VGND VGND VPWR VPWR _15283_/X sky130_fd_sc_hd__and3_4
XFILLER_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17378__A _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12494_/X VGND VGND VPWR VPWR _12495_/Y sky130_fd_sc_hd__inv_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _16008_/Y _24408_/Q _16008_/Y _24408_/Q VGND VGND VPWR VPWR _17022_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14234_ _14227_/Y _14233_/X _13844_/X _14233_/X VGND VGND VPWR VPWR _14234_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14165_ _25221_/Q _14109_/B _25221_/Q _14109_/B VGND VGND VPWR VPWR _14165_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13116_ _12342_/Y _13115_/X VGND VGND VPWR VPWR _13121_/A sky130_fd_sc_hd__or2_4
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21628__A _14761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14096_ _13994_/A _14090_/X _14087_/X _14027_/D _14093_/X VGND VGND VPWR VPWR _25235_/D
+ sky130_fd_sc_hd__a32o_4
X_18973_ _18973_/A VGND VGND VPWR VPWR _18973_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13489__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13047_ _13044_/A _13039_/B _13046_/X VGND VGND VPWR VPWR _13047_/X sky130_fd_sc_hd__and3_4
X_17924_ _15923_/B _17924_/B VGND VGND VPWR VPWR _17924_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15626__A _15626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19613__B1 _19612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17855_ _17896_/A VGND VGND VPWR VPWR _17881_/A sky130_fd_sc_hd__buf_2
XFILLER_121_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17263__D _17262_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16806_ _16805_/X VGND VGND VPWR VPWR _16806_/X sky130_fd_sc_hd__buf_2
X_17786_ _17788_/B VGND VGND VPWR VPWR _17787_/B sky130_fd_sc_hd__inv_2
X_14998_ _15243_/A _16770_/A _15243_/A _16770_/A VGND VGND VPWR VPWR _14998_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19525_ _21199_/B _19520_/X _19501_/X _19507_/Y VGND VGND VPWR VPWR _23717_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16737_ _16468_/A _16382_/B VGND VGND VPWR VPWR _16737_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13949_ _13949_/A VGND VGND VPWR VPWR _13949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16457__A _18515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21723__B2 _21535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_191_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _23395_/CLK sky130_fd_sc_hd__clkbuf_1
X_19456_ _18214_/B VGND VGND VPWR VPWR _19456_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16668_ _16666_/Y _16667_/X _16309_/X _16667_/X VGND VGND VPWR VPWR _16668_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18407_ _24184_/Q VGND VGND VPWR VPWR _18534_/A sky130_fd_sc_hd__inv_2
XFILLER_201_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_48_0_HCLK clkbuf_7_24_0_HCLK/X VGND VGND VPWR VPWR _25292_/CLK sky130_fd_sc_hd__clkbuf_1
X_15619_ _15618_/Y _15614_/X _11827_/X _15614_/X VGND VGND VPWR VPWR _24909_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22279__A2 _22259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19387_ _18206_/B VGND VGND VPWR VPWR _19387_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16599_ _24533_/Q VGND VGND VPWR VPWR _16599_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_29_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24590__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _18938_/A _18333_/X _19815_/A VGND VGND VPWR VPWR _18338_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_187_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18269_ _18268_/X _20405_/A VGND VGND VPWR VPWR _18269_/X sky130_fd_sc_hd__or2_4
XANTENNA__16192__A _16192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16902__B2 _16910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20300_ _20300_/A VGND VGND VPWR VPWR _22344_/B sky130_fd_sc_hd__inv_2
XANTENNA__21239__B1 _21229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21280_ _21280_/A VGND VGND VPWR VPWR _21386_/B sky130_fd_sc_hd__buf_2
X_20231_ _20230_/Y _20226_/X _20146_/X _20213_/Y VGND VGND VPWR VPWR _20231_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15469__A1 _14289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__B _21104_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20162_ _23495_/Q VGND VGND VPWR VPWR _21647_/B sky130_fd_sc_hd__inv_2
XANTENNA__21538__A _21129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20093_ _20093_/A VGND VGND VPWR VPWR _20093_/X sky130_fd_sc_hd__buf_2
X_24970_ _24975_/CLK _24970_/D HRESETn VGND VGND VPWR VPWR _13910_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22203__A2 _22425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19604__B1 _19418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19008__A _19148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16418__B1 _16417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23921_ _25491_/CLK _23921_/D VGND VGND VPWR VPWR _23921_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19080__B2 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17751__A _17751_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23852_ _23885_/CLK _23852_/D VGND VGND VPWR VPWR _19141_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22803_ _16689_/Y _22890_/B VGND VGND VPWR VPWR _22803_/X sky130_fd_sc_hd__and2_4
XFILLER_226_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23783_ _24252_/CLK _23783_/D VGND VGND VPWR VPWR _23783_/Q sky130_fd_sc_hd__dfxtp_4
X_20995_ _20996_/A _20995_/B _20996_/C VGND VGND VPWR VPWR _23943_/D sky130_fd_sc_hd__and3_4
XANTENNA__16367__A _24620_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17918__B1 _22003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22911__B1 _24844_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25522_ _25520_/CLK _11907_/X HRESETn VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__dfrtp_4
X_22734_ _22733_/X VGND VGND VPWR VPWR _22734_/Y sky130_fd_sc_hd__inv_2
XFILLER_214_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24678__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20168__A2_N _20163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25453_ _25454_/CLK _25453_/D HRESETn VGND VGND VPWR VPWR _12257_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24607__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22665_ _22665_/A _22662_/B VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__or2_4
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24404_ _24952_/CLK _17085_/Y HRESETn VGND VGND VPWR VPWR _24404_/Q sky130_fd_sc_hd__dfrtp_4
X_21616_ _21648_/A _19270_/Y VGND VGND VPWR VPWR _21616_/X sky130_fd_sc_hd__or2_4
XFILLER_187_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25384_ _25402_/CLK _25384_/D HRESETn VGND VGND VPWR VPWR _12955_/A sky130_fd_sc_hd__dfrtp_4
X_22596_ _22523_/X _22594_/X _21968_/X _22595_/X VGND VGND VPWR VPWR _22596_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24337_/CLK _24335_/D HRESETn VGND VGND VPWR VPWR _24335_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23219__A1 _24579_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21547_ _21126_/B VGND VGND VPWR VPWR _21547_/X sky130_fd_sc_hd__buf_2
XFILLER_194_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12280_ _12274_/X _12280_/B _12280_/C _12279_/X VGND VGND VPWR VPWR _12281_/D sky130_fd_sc_hd__or4_4
X_24266_ _24715_/CLK _17890_/X HRESETn VGND VGND VPWR VPWR _24266_/Q sky130_fd_sc_hd__dfrtp_4
X_21478_ _21482_/A _21478_/B _21477_/X VGND VGND VPWR VPWR _21478_/X sky130_fd_sc_hd__and3_4
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23217_ _23249_/A _23216_/Y VGND VGND VPWR VPWR _23217_/Y sky130_fd_sc_hd__nor2_4
X_20429_ _13316_/B VGND VGND VPWR VPWR _20429_/Y sky130_fd_sc_hd__inv_2
X_24197_ _24196_/CLK _24197_/D HRESETn VGND VGND VPWR VPWR _18393_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21650__B1 _14758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23148_ _23148_/A VGND VGND VPWR VPWR _23148_/X sky130_fd_sc_hd__buf_2
XANTENNA__21448__A _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15970_ HWDATA[18] VGND VGND VPWR VPWR _15970_/X sky130_fd_sc_hd__buf_2
X_23079_ _23013_/A _23076_/X _23079_/C VGND VGND VPWR VPWR _23079_/X sky130_fd_sc_hd__and3_4
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21167__B _21172_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14921_ _14921_/A VGND VGND VPWR VPWR _14921_/X sky130_fd_sc_hd__buf_2
XFILLER_209_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13891__B1 _23444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17640_ _17579_/A _17637_/X VGND VGND VPWR VPWR _17640_/X sky130_fd_sc_hd__or2_4
XFILLER_208_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14852_ _14852_/A VGND VGND VPWR VPWR _14852_/X sky130_fd_sc_hd__buf_2
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13803_ _21384_/B VGND VGND VPWR VPWR _13804_/D sky130_fd_sc_hd__buf_2
X_14783_ _14783_/A _14785_/A _14785_/B VGND VGND VPWR VPWR _14783_/X sky130_fd_sc_hd__and3_4
X_17571_ _24319_/Q VGND VGND VPWR VPWR _17571_/Y sky130_fd_sc_hd__inv_2
X_11995_ _11663_/A _11992_/X _11987_/Y _11994_/Y VGND VGND VPWR VPWR _25502_/D sky130_fd_sc_hd__o22a_4
XFILLER_17_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21705__A1 _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19310_ _19307_/Y _19302_/X _19308_/X _19309_/X VGND VGND VPWR VPWR _23794_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_217_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_201_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24189_/CLK sky130_fd_sc_hd__clkbuf_1
X_13734_ _13693_/A _13692_/X VGND VGND VPWR VPWR _13734_/Y sky130_fd_sc_hd__nand2_4
X_16522_ _16522_/A VGND VGND VPWR VPWR _16522_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_7_0_HCLK clkbuf_8_6_0_HCLK/A VGND VGND VPWR VPWR _24217_/CLK sky130_fd_sc_hd__clkbuf_1
X_19241_ _19249_/A VGND VGND VPWR VPWR _19241_/X sky130_fd_sc_hd__buf_2
XFILLER_220_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21911__A _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13665_ _24051_/Q _13664_/X VGND VGND VPWR VPWR _13666_/B sky130_fd_sc_hd__or2_4
X_16453_ _15134_/Y _16384_/A _16276_/X _16384_/A VGND VGND VPWR VPWR _24586_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15935__A2 _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22726__B _21877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12616_ _12616_/A _12616_/B VGND VGND VPWR VPWR _12629_/C sky130_fd_sc_hd__or2_4
X_15404_ _15407_/A _15407_/B VGND VGND VPWR VPWR _15408_/B sky130_fd_sc_hd__or2_4
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16384_ _16384_/A VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__buf_2
X_19172_ _19171_/Y _19168_/X _19148_/X _19168_/X VGND VGND VPWR VPWR _19172_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13596_ _13590_/X _13596_/B _13594_/X _13595_/X VGND VGND VPWR VPWR _13596_/X sky130_fd_sc_hd__or4_4
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15335_ _15302_/Y _15334_/X _15324_/X _15331_/B VGND VGND VPWR VPWR _15336_/A sky130_fd_sc_hd__a211o_4
X_18123_ _18234_/A _18119_/X _18123_/C VGND VGND VPWR VPWR _18123_/X sky130_fd_sc_hd__or3_4
X_12547_ _25430_/Q VGND VGND VPWR VPWR _12616_/B sky130_fd_sc_hd__inv_2
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15266_ _15260_/C _15265_/X _14996_/X _15261_/Y VGND VGND VPWR VPWR _15266_/X sky130_fd_sc_hd__a211o_4
X_18054_ _18127_/A _18052_/X _18054_/C VGND VGND VPWR VPWR _18054_/X sky130_fd_sc_hd__and3_4
X_12478_ _12291_/D _12478_/B VGND VGND VPWR VPWR _12479_/B sky130_fd_sc_hd__or2_4
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22969__B1 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _20525_/B _14208_/X _13806_/X _14210_/X VGND VGND VPWR VPWR _14217_/X sky130_fd_sc_hd__a2bb2o_4
X_17005_ _16053_/Y _24390_/Q _16053_/Y _24390_/Q VGND VGND VPWR VPWR _17005_/X sky130_fd_sc_hd__a2bb2o_4
X_15197_ _15068_/X _15197_/B _15197_/C VGND VGND VPWR VPWR _15197_/X sky130_fd_sc_hd__and3_4
XFILLER_153_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14148_ _25226_/Q _14125_/X _25226_/Q _14125_/X VGND VGND VPWR VPWR _14149_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14079_ _14060_/A _14040_/Y VGND VGND VPWR VPWR _14079_/X sky130_fd_sc_hd__or2_4
X_18956_ _23917_/Q VGND VGND VPWR VPWR _18956_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17907_ _17907_/A _17907_/B VGND VGND VPWR VPWR _17907_/X sky130_fd_sc_hd__and2_4
XFILLER_140_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18887_ _18887_/A _18887_/B VGND VGND VPWR VPWR _18888_/B sky130_fd_sc_hd__or2_4
X_17838_ _17768_/D _17820_/B _17790_/X _17836_/B VGND VGND VPWR VPWR _17839_/A sky130_fd_sc_hd__a211o_4
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17769_ _17762_/Y _17763_/Y _17766_/X _17769_/D VGND VGND VPWR VPWR _17770_/B sky130_fd_sc_hd__or4_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _19507_/Y VGND VGND VPWR VPWR _19508_/X sky130_fd_sc_hd__buf_2
XFILLER_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13604__A _19548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24771__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20780_ _20779_/X VGND VGND VPWR VPWR _20780_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17376__A1 _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22917__A _24636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21821__A _21687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24700__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19439_ _19032_/A VGND VGND VPWR VPWR _19439_/X sky130_fd_sc_hd__buf_2
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20380__B1 _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22450_ _22732_/A _22448_/X _21456_/X _22449_/X VGND VGND VPWR VPWR _22450_/X sky130_fd_sc_hd__o22a_4
XFILLER_210_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21401_ _21412_/A _21399_/X _21401_/C VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__and3_4
X_22381_ _22385_/A _18912_/Y VGND VGND VPWR VPWR _22383_/B sky130_fd_sc_hd__or2_4
XANTENNA__14435__A _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24120_ _23954_/CLK _24120_/D HRESETn VGND VGND VPWR VPWR _24120_/Q sky130_fd_sc_hd__dfrtp_4
X_21332_ _21332_/A _21173_/C VGND VGND VPWR VPWR _21332_/X sky130_fd_sc_hd__or2_4
XFILLER_129_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24051_ _24488_/CLK _20853_/Y HRESETn VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfrtp_4
X_21263_ _21263_/A _20188_/Y VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__or2_4
XFILLER_237_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19825__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23002_ _16677_/Y _23177_/B VGND VGND VPWR VPWR _23002_/X sky130_fd_sc_hd__and2_4
X_20214_ _20213_/Y VGND VGND VPWR VPWR _20214_/X sky130_fd_sc_hd__buf_2
XFILLER_190_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21194_ _21207_/A _21194_/B VGND VGND VPWR VPWR _21194_/X sky130_fd_sc_hd__or2_4
XFILLER_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20145_ _20145_/A VGND VGND VPWR VPWR _20145_/Y sky130_fd_sc_hd__inv_2
X_24953_ _24952_/CLK _15502_/X HRESETn VGND VGND VPWR VPWR _12061_/A sky130_fd_sc_hd__dfrtp_4
X_20076_ _20076_/A VGND VGND VPWR VPWR _21271_/B sky130_fd_sc_hd__inv_2
XFILLER_246_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20900__A _20836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23904_ _23885_/CLK _18993_/X VGND VGND VPWR VPWR _23904_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24859__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24884_ _24889_/CLK _15736_/X HRESETn VGND VGND VPWR VPWR _24884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21715__B _22897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23835_ _23850_/CLK _23835_/D VGND VGND VPWR VPWR _19193_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16097__A _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ HWDATA[23] VGND VGND VPWR VPWR _11780_/X sky130_fd_sc_hd__buf_2
X_23766_ _23768_/CLK _23766_/D VGND VGND VPWR VPWR _19385_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20978_ _24113_/Q _12172_/B VGND VGND VPWR VPWR _20978_/Y sky130_fd_sc_hd__nor2_4
XFILLER_26_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21163__A2 _14229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22717_ _16512_/A _21855_/B _21096_/X VGND VGND VPWR VPWR _22717_/X sky130_fd_sc_hd__and3_4
X_25505_ _25507_/CLK _11980_/Y HRESETn VGND VGND VPWR VPWR _25505_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23697_ _23441_/CLK _19583_/X VGND VGND VPWR VPWR _19582_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_186_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16825__A _16810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13450_ _13450_/A _18979_/A VGND VGND VPWR VPWR _13451_/C sky130_fd_sc_hd__or2_4
X_25436_ _25419_/CLK _25436_/D HRESETn VGND VGND VPWR VPWR _12601_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_31_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24732_/CLK sky130_fd_sc_hd__clkbuf_1
X_22648_ _21082_/A _22645_/X _21116_/X _22647_/X VGND VGND VPWR VPWR _22648_/Y sky130_fd_sc_hd__a22oi_4
X_12401_ _12225_/Y _12401_/B _12401_/C VGND VGND VPWR VPWR _12401_/X sky130_fd_sc_hd__or3_4
XFILLER_167_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_94_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _24889_/CLK sky130_fd_sc_hd__clkbuf_1
X_13381_ _13413_/A _13381_/B VGND VGND VPWR VPWR _13381_/X sky130_fd_sc_hd__or2_4
X_25367_ _25365_/CLK _25367_/D HRESETn VGND VGND VPWR VPWR _12306_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22579_ _21123_/A _22577_/X _22121_/X _22578_/X VGND VGND VPWR VPWR _22580_/B sky130_fd_sc_hd__o22a_4
XFILLER_194_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17359__C _17359_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15120_ _24990_/Q VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__inv_2
X_12332_ _25347_/Q VGND VGND VPWR VPWR _12332_/Y sky130_fd_sc_hd__inv_2
X_24318_ _24327_/CLK _24318_/D HRESETn VGND VGND VPWR VPWR _17553_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21871__B1 _21121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25298_ _24406_/CLK _25298_/D HRESETn VGND VGND VPWR VPWR _13702_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15051_ _15051_/A VGND VGND VPWR VPWR _15051_/Y sky130_fd_sc_hd__inv_2
X_12263_ _25442_/Q VGND VGND VPWR VPWR _12263_/Y sky130_fd_sc_hd__inv_2
X_24249_ _24252_/CLK _24249_/D HRESETn VGND VGND VPWR VPWR _24249_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15550__B1 HADDR[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22415__A2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14002_ _14062_/A _14042_/B _14032_/A _14001_/X VGND VGND VPWR VPWR _14003_/A sky130_fd_sc_hd__or4_4
XFILLER_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12194_ _12428_/A _24778_/Q _12428_/A _24778_/Q VGND VGND VPWR VPWR _12195_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18810_ _18810_/A _18810_/B VGND VGND VPWR VPWR _18810_/X sky130_fd_sc_hd__or2_4
X_19790_ _16866_/X VGND VGND VPWR VPWR _19790_/X sky130_fd_sc_hd__buf_2
X_18741_ _18683_/B _18735_/B _18740_/X _18736_/Y VGND VGND VPWR VPWR _18742_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15953_ _15947_/A VGND VGND VPWR VPWR _15953_/X sky130_fd_sc_hd__buf_2
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14904_ _15206_/A _24444_/Q _14902_/Y _24444_/Q VGND VGND VPWR VPWR _14904_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17391__A _17391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18672_ _16617_/Y _24137_/Q _16625_/Y _24134_/Q VGND VGND VPWR VPWR _18672_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15884_ _12781_/Y _15880_/X _11776_/X _15880_/X VGND VGND VPWR VPWR _15884_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16802__B1 _16729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17623_ _17520_/Y _17626_/B VGND VGND VPWR VPWR _17627_/B sky130_fd_sc_hd__or2_4
XANTENNA__24529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14835_ _14835_/A VGND VGND VPWR VPWR _14840_/A sky130_fd_sc_hd__buf_2
XFILLER_205_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ _25547_/Q _17553_/Y _11789_/Y _24316_/Q VGND VGND VPWR VPWR _17554_/X sky130_fd_sc_hd__a2bb2o_4
X_11978_ _25505_/Q VGND VGND VPWR VPWR _11978_/Y sky130_fd_sc_hd__inv_2
X_14766_ _14765_/X VGND VGND VPWR VPWR _14766_/X sky130_fd_sc_hd__buf_2
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16505_ _16504_/Y _16500_/X _16419_/X _16500_/X VGND VGND VPWR VPWR _16505_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _11666_/Y _13700_/B VGND VGND VPWR VPWR _13717_/Y sky130_fd_sc_hd__nand2_4
X_14697_ _21263_/A VGND VGND VPWR VPWR _21914_/A sky130_fd_sc_hd__buf_2
X_17485_ _17484_/A VGND VGND VPWR VPWR _17485_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19224_ _18168_/B VGND VGND VPWR VPWR _19224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16436_ _16434_/Y _16435_/X _16252_/X _16435_/X VGND VGND VPWR VPWR _24596_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ _13547_/Y _13642_/X _13647_/X VGND VGND VPWR VPWR _25307_/D sky130_fd_sc_hd__a21oi_4
XANTENNA__23300__B1 _24293_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19155_ _19154_/Y _19152_/X _19085_/X _19152_/X VGND VGND VPWR VPWR _19155_/X sky130_fd_sc_hd__a2bb2o_4
X_13579_ _13577_/A VGND VGND VPWR VPWR _14590_/A sky130_fd_sc_hd__inv_2
X_16367_ _24620_/Q VGND VGND VPWR VPWR _16367_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_2_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18106_ _18138_/A _18106_/B _18105_/X VGND VGND VPWR VPWR _18107_/C sky130_fd_sc_hd__or3_4
XFILLER_117_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16869__B1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15318_ _15302_/Y _15340_/A _15318_/C _15337_/B VGND VGND VPWR VPWR _15318_/X sky130_fd_sc_hd__or4_4
X_16298_ _16325_/A VGND VGND VPWR VPWR _16298_/X sky130_fd_sc_hd__buf_2
X_19086_ _19084_/Y _19082_/X _19085_/X _19082_/X VGND VGND VPWR VPWR _23873_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22472__A _22472_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17530__A1 _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18037_ _18037_/A _18037_/B _18036_/X VGND VGND VPWR VPWR _18037_/X sky130_fd_sc_hd__and3_4
X_15249_ _15249_/A VGND VGND VPWR VPWR _15249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15541__B1 HADDR[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21088__A _22968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22811__C1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19988_ _19988_/A VGND VGND VPWR VPWR _19988_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14647__A2 _13610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18939_ _18938_/X VGND VGND VPWR VPWR _18952_/A sky130_fd_sc_hd__inv_2
X_21950_ _21945_/X _21949_/X _18306_/A VGND VGND VPWR VPWR _21950_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16934__A2_N _17832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20901_ _13672_/X VGND VGND VPWR VPWR _20907_/B sky130_fd_sc_hd__buf_2
XFILLER_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21881_ _21430_/X VGND VGND VPWR VPWR _21881_/X sky130_fd_sc_hd__buf_2
XFILLER_227_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18609__A1_N _16617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23620_ _23916_/CLK _19818_/X VGND VGND VPWR VPWR _23620_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _20881_/A VGND VGND VPWR VPWR _20854_/A sky130_fd_sc_hd__buf_2
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21551__A _21436_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _23534_/CLK _23551_/D VGND VGND VPWR VPWR _23551_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20763_ _20768_/B VGND VGND VPWR VPWR _20763_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20353__B1 _20243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22502_ _22502_/A _22662_/B VGND VGND VPWR VPWR _22502_/X sky130_fd_sc_hd__or2_4
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22134__A2_N _22176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _24684_/CLK _23482_/D VGND VGND VPWR VPWR _23482_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20694_ _20694_/A VGND VGND VPWR VPWR _20716_/A sky130_fd_sc_hd__buf_2
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25221_ _25223_/CLK _14167_/X HRESETn VGND VGND VPWR VPWR _25221_/Q sky130_fd_sc_hd__dfrtp_4
X_22433_ _25380_/Q _22306_/X _22432_/X VGND VGND VPWR VPWR _22433_/X sky130_fd_sc_hd__a21o_4
XANTENNA__15780__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25152_ _25154_/CLK _25152_/D HRESETn VGND VGND VPWR VPWR _25152_/Q sky130_fd_sc_hd__dfrtp_4
X_22364_ _21473_/A _22364_/B VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__or2_4
XFILLER_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24103_ _25188_/CLK _24103_/D HRESETn VGND VGND VPWR VPWR _20971_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21315_ _21332_/A VGND VGND VPWR VPWR _22577_/B sky130_fd_sc_hd__buf_2
X_25083_ _23885_/CLK _14651_/X HRESETn VGND VGND VPWR VPWR _25083_/Q sky130_fd_sc_hd__dfrtp_4
X_22295_ _21101_/X VGND VGND VPWR VPWR _23299_/A sky130_fd_sc_hd__buf_2
XANTENNA__16380__A _14199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24034_ _24495_/CLK _20783_/Y HRESETn VGND VGND VPWR VPWR _24034_/Q sky130_fd_sc_hd__dfrtp_4
X_21246_ _21246_/A VGND VGND VPWR VPWR _21638_/A sky130_fd_sc_hd__buf_2
XANTENNA__19274__B2 _19271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21177_ _21177_/A _21177_/B _21177_/C VGND VGND VPWR VPWR _21226_/C sky130_fd_sc_hd__and3_4
XFILLER_132_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20128_ _20128_/A VGND VGND VPWR VPWR _20129_/A sky130_fd_sc_hd__buf_2
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12950_ _12854_/X _12988_/B VGND VGND VPWR VPWR _12950_/X sky130_fd_sc_hd__or2_4
XANTENNA__24693__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _20059_/A VGND VGND VPWR VPWR _20059_/Y sky130_fd_sc_hd__inv_2
X_24936_ _24937_/CLK _24936_/D HRESETn VGND VGND VPWR VPWR _21135_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_86_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11901_ _11901_/A _11898_/B VGND VGND VPWR VPWR _11902_/A sky130_fd_sc_hd__or2_4
XANTENNA__24622__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12881_ _12790_/Y _12878_/X VGND VGND VPWR VPWR _12881_/X sky130_fd_sc_hd__or2_4
XFILLER_245_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24867_ _24867_/CLK _24867_/D HRESETn VGND VGND VPWR VPWR _24867_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11829_/Y _11825_/X _11831_/X _11825_/X VGND VGND VPWR VPWR _25535_/D sky130_fd_sc_hd__a2bb2o_4
X_14620_ _14570_/B _14619_/X _14566_/X _14611_/X _13561_/A VGND VGND VPWR VPWR _25089_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _23454_/CLK _19242_/X VGND VGND VPWR VPWR _13274_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24798_ _24781_/CLK _24798_/D HRESETn VGND VGND VPWR VPWR _24798_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14271__B1 _13846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14544_/Y _14082_/B _20461_/C VGND VGND VPWR VPWR _14551_/X sky130_fd_sc_hd__o21a_4
XFILLER_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ HWDATA[28] VGND VGND VPWR VPWR _11763_/X sky130_fd_sc_hd__buf_2
X_23749_ _23735_/CLK _23749_/D VGND VGND VPWR VPWR _18213_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13502_/A VGND VGND VPWR VPWR _13502_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14481_/Y _14475_/X _14409_/X _14468_/A VGND VGND VPWR VPWR _14482_/X sky130_fd_sc_hd__a2bb2o_4
X_17270_ _17203_/Y _17243_/X _17270_/C _17283_/B VGND VGND VPWR VPWR _17271_/A sky130_fd_sc_hd__or4_4
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11694_/A VGND VGND VPWR VPWR _13697_/A sky130_fd_sc_hd__inv_2
XFILLER_41_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13433_ _13369_/A _13433_/B VGND VGND VPWR VPWR _13434_/C sky130_fd_sc_hd__or2_4
X_16221_ _24673_/Q VGND VGND VPWR VPWR _16221_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25419_ _25419_/CLK _25419_/D HRESETn VGND VGND VPWR VPWR _25419_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15771__B1 _15632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16152_ _22502_/A VGND VGND VPWR VPWR _16152_/Y sky130_fd_sc_hd__inv_2
X_13364_ _13249_/A _23792_/Q VGND VGND VPWR VPWR _13366_/B sky130_fd_sc_hd__or2_4
XFILLER_6_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12315_ _25366_/Q VGND VGND VPWR VPWR _13026_/A sky130_fd_sc_hd__inv_2
X_15103_ _15103_/A _15097_/X _15100_/X _15102_/X VGND VGND VPWR VPWR _15103_/X sky130_fd_sc_hd__or4_4
X_16083_ _16082_/Y _16005_/X _15848_/X _16005_/X VGND VGND VPWR VPWR _16083_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17386__A _17389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15523__B1 HADDR[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13295_ _13428_/A _13295_/B VGND VGND VPWR VPWR _13295_/X sky130_fd_sc_hd__or2_4
XFILLER_6_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16290__A _16290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15034_ _24472_/Q VGND VGND VPWR VPWR _15034_/Y sky130_fd_sc_hd__inv_2
X_19911_ _19909_/Y _19905_/X _19632_/X _19910_/X VGND VGND VPWR VPWR _19911_/X sky130_fd_sc_hd__a2bb2o_4
X_12246_ _12246_/A VGND VGND VPWR VPWR _12247_/A sky130_fd_sc_hd__inv_2
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21072__A1 _24719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19842_ _22230_/B _19839_/X _19793_/X _19839_/X VGND VGND VPWR VPWR _23611_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13419__A _13451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12177_ _12177_/A VGND VGND VPWR VPWR _12177_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21636__A _22090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19773_ _19765_/Y VGND VGND VPWR VPWR _19773_/X sky130_fd_sc_hd__buf_2
XFILLER_228_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16985_ _24402_/Q VGND VGND VPWR VPWR _17088_/A sky130_fd_sc_hd__inv_2
XANTENNA__13837__B1 _11827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18724_ _18710_/A _18702_/X VGND VGND VPWR VPWR _18727_/B sky130_fd_sc_hd__or2_4
X_15936_ _15683_/X _15934_/B VGND VGND VPWR VPWR _15936_/X sky130_fd_sc_hd__or2_4
XFILLER_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18655_ _16574_/Y _18744_/A _16574_/Y _24154_/Q VGND VGND VPWR VPWR _18659_/B sky130_fd_sc_hd__a2bb2o_4
X_15867_ _15866_/X VGND VGND VPWR VPWR _23053_/A sky130_fd_sc_hd__buf_2
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18945__A _18952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17606_ _17525_/A _17606_/B VGND VGND VPWR VPWR _17608_/B sky130_fd_sc_hd__or2_4
XFILLER_91_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13154__A _13153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14818_ _14835_/A VGND VGND VPWR VPWR _14837_/A sky130_fd_sc_hd__inv_2
X_18586_ _18569_/X _18586_/B _18598_/C VGND VGND VPWR VPWR _18586_/X sky130_fd_sc_hd__and3_4
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15798_ _15715_/X VGND VGND VPWR VPWR _21043_/A sky130_fd_sc_hd__buf_2
XFILLER_212_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22467__A _16284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17537_ _24297_/Q VGND VGND VPWR VPWR _17537_/Y sky130_fd_sc_hd__inv_2
X_14749_ _22056_/A _14749_/B VGND VGND VPWR VPWR _14749_/X sky130_fd_sc_hd__or2_4
XANTENNA__12812__B2 _22726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17468_ _17466_/A _17465_/X _18347_/A _17467_/Y VGND VGND VPWR VPWR _17471_/A sky130_fd_sc_hd__o22a_4
X_19207_ _18231_/B VGND VGND VPWR VPWR _19207_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16419_ HWDATA[17] VGND VGND VPWR VPWR _16419_/X sky130_fd_sc_hd__buf_2
XFILLER_220_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15762__B1 _24871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17399_ _17399_/A _17399_/B VGND VGND VPWR VPWR _17399_/X sky130_fd_sc_hd__or2_4
X_19138_ _23853_/Q VGND VGND VPWR VPWR _19138_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14317__A1 MSO_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19069_ _19067_/Y _19068_/X _18975_/X _19068_/X VGND VGND VPWR VPWR _19069_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15514__B1 HADDR[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14713__A _14713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21100_ _24825_/Q _21085_/X _21042_/X _21099_/X VGND VGND VPWR VPWR _21100_/X sky130_fd_sc_hd__a211o_4
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22080_ _22085_/A _22080_/B VGND VGND VPWR VPWR _22080_/X sky130_fd_sc_hd__or2_4
XANTENNA__22930__A _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21031_ _21031_/A VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__buf_2
XANTENNA__12233__A _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15544__A _15544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22982_ _22982_/A _23158_/B VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__or2_4
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21933_ _21938_/A _21933_/B VGND VGND VPWR VPWR _21933_/X sky130_fd_sc_hd__or2_4
X_24721_ _24726_/CLK _16085_/X HRESETn VGND VGND VPWR VPWR _24721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24652_ _24169_/CLK _24652_/D HRESETn VGND VGND VPWR VPWR _16278_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23107__A3 _22291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21864_ _12122_/Y _12107_/X _18386_/Y _12080_/X VGND VGND VPWR VPWR _21864_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23603_ _25068_/CLK _19865_/X VGND VGND VPWR VPWR _23603_/Q sky130_fd_sc_hd__dfxtp_4
X_20815_ _23213_/A _20716_/A _20788_/A _20814_/Y VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__o22a_4
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24583_ _24562_/CLK _24583_/D HRESETn VGND VGND VPWR VPWR _16466_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21795_ _21777_/X _21794_/X _22400_/A VGND VGND VPWR VPWR _21795_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12803__B2 _22139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23534_/CLK _23534_/D VGND VGND VPWR VPWR _20053_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_168_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20746_ _20746_/A VGND VGND VPWR VPWR _20746_/Y sky130_fd_sc_hd__inv_2
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23466_/CLK _23465_/D VGND VGND VPWR VPWR _23465_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15753__B1 _24875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20677_ _14235_/Y _20622_/Y _20637_/A _20676_/Y VGND VGND VPWR VPWR _20677_/X sky130_fd_sc_hd__a211o_4
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25204_ _25204_/CLK _14239_/X HRESETn VGND VGND VPWR VPWR _20672_/A sky130_fd_sc_hd__dfstp_4
XFILLER_149_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22416_ _24270_/Q _21113_/X _21711_/A VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__o21a_4
X_23396_ _24206_/CLK _20418_/X VGND VGND VPWR VPWR _21218_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_192_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_105_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24015_/CLK sky130_fd_sc_hd__clkbuf_1
X_25135_ _25137_/CLK _25135_/D HRESETn VGND VGND VPWR VPWR _25135_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__23001__A _22999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22347_ _21938_/A _22347_/B VGND VGND VPWR VPWR _22348_/C sky130_fd_sc_hd__or2_4
XANTENNA__15505__B1 HADDR[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_168_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23830_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12100_ _12099_/Y _12095_/X _11876_/X _12083_/A VGND VGND VPWR VPWR _12100_/X sky130_fd_sc_hd__a2bb2o_4
X_13080_ _13021_/C _13006_/C VGND VGND VPWR VPWR _13080_/X sky130_fd_sc_hd__or2_4
X_25066_ _25066_/CLK _25066_/D HRESETn VGND VGND VPWR VPWR _21240_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22278_ _11670_/Y _21513_/X _21519_/X VGND VGND VPWR VPWR _22278_/X sky130_fd_sc_hd__a21o_4
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14342__B _14342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12031_ _12029_/A _12030_/A _12029_/Y _12030_/Y VGND VGND VPWR VPWR _12035_/C sky130_fd_sc_hd__o22a_4
X_24017_ _24485_/CLK _20707_/Y HRESETn VGND VGND VPWR VPWR _24017_/Q sky130_fd_sc_hd__dfrtp_4
X_21229_ _22808_/A VGND VGND VPWR VPWR _21229_/X sky130_fd_sc_hd__buf_2
XANTENNA__24874__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21456__A _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24803__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16770_ _16770_/A VGND VGND VPWR VPWR _16770_/Y sky130_fd_sc_hd__inv_2
X_13982_ _13982_/A _13982_/B VGND VGND VPWR VPWR _13982_/X sky130_fd_sc_hd__or2_4
XANTENNA__21357__A2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22554__A1 _17359_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15721_ _15557_/X _15714_/X _15562_/X _24891_/Q _15720_/X VGND VGND VPWR VPWR _15721_/X
+ sky130_fd_sc_hd__a32o_4
X_12933_ _12912_/B _12911_/X VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__or2_4
X_24919_ _24923_/CLK _15595_/X HRESETn VGND VGND VPWR VPWR _15594_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_206_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18440_ _16217_/Y _24186_/Q _16217_/Y _24186_/Q VGND VGND VPWR VPWR _18443_/B sky130_fd_sc_hd__a2bb2o_4
X_15652_ _15651_/X VGND VGND VPWR VPWR _15652_/Y sky130_fd_sc_hd__inv_2
X_12864_ _12864_/A _12863_/X VGND VGND VPWR VPWR _12872_/A sky130_fd_sc_hd__or2_4
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14603_/A _14575_/X VGND VGND VPWR VPWR _14603_/Y sky130_fd_sc_hd__nand2_4
XFILLER_221_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11815_ _11811_/Y _11804_/X _11813_/X _11814_/X VGND VGND VPWR VPWR _25539_/D sky130_fd_sc_hd__a2bb2o_4
X_18371_ _18363_/X _18370_/Y _24206_/Q _18362_/Y VGND VGND VPWR VPWR _24206_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12793_/A _22490_/A _12855_/A _12794_/Y VGND VGND VPWR VPWR _12799_/C sky130_fd_sc_hd__o22a_4
X_15583_ _15583_/A VGND VGND VPWR VPWR _15583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22857__A2 _22841_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15992__B1 _24757_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16285__A _16284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17322_/A _17322_/B VGND VGND VPWR VPWR _17323_/C sky130_fd_sc_hd__or2_4
XFILLER_187_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _22575_/A VGND VGND VPWR VPWR _11747_/A sky130_fd_sc_hd__buf_2
X_14534_ _14530_/X _14533_/X _14492_/A _14526_/X VGND VGND VPWR VPWR _25111_/D sky130_fd_sc_hd__o22a_4
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _17253_/A VGND VGND VPWR VPWR _17253_/Y sky130_fd_sc_hd__inv_2
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11676_/Y _24238_/Q _11676_/Y _24238_/Q VGND VGND VPWR VPWR _11677_/X sky130_fd_sc_hd__a2bb2o_4
X_14465_ _14465_/A VGND VGND VPWR VPWR _14465_/Y sky130_fd_sc_hd__inv_2
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12318__A _24852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16204_ _16201_/Y _16197_/X _15948_/X _16203_/X VGND VGND VPWR VPWR _16204_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13416_ _13416_/A _13416_/B _13415_/X VGND VGND VPWR VPWR _13424_/B sky130_fd_sc_hd__or3_4
Xclkbuf_7_64_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_64_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14396_ _14395_/Y _14391_/X _13846_/X _14393_/X VGND VGND VPWR VPWR _14396_/X sky130_fd_sc_hd__a2bb2o_4
X_17184_ _17184_/A VGND VGND VPWR VPWR _17359_/C sky130_fd_sc_hd__buf_2
XANTENNA__17828__B _17832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13347_ _13411_/A _19130_/A VGND VGND VPWR VPWR _13348_/C sky130_fd_sc_hd__or2_4
X_16135_ _16096_/X VGND VGND VPWR VPWR _16162_/A sky130_fd_sc_hd__buf_2
XANTENNA__15629__A _14420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18005__A _18102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13278_ _13385_/A _13278_/B VGND VGND VPWR VPWR _13278_/X sky130_fd_sc_hd__or2_4
X_16066_ _14420_/A VGND VGND VPWR VPWR _16066_/X sky130_fd_sc_hd__buf_2
X_12229_ _12228_/Y VGND VGND VPWR VPWR _12229_/X sky130_fd_sc_hd__buf_2
X_15017_ _15017_/A VGND VGND VPWR VPWR _15017_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18997__B1 _18908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19825_ _19824_/Y _19822_/X _19728_/X _19822_/X VGND VGND VPWR VPWR _19825_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19756_ _19742_/Y VGND VGND VPWR VPWR _19756_/X sky130_fd_sc_hd__buf_2
X_16968_ _15999_/Y _17062_/A _15999_/Y _17062_/A VGND VGND VPWR VPWR _16972_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18707_ _18606_/X _18708_/B VGND VGND VPWR VPWR _18709_/B sky130_fd_sc_hd__or2_4
X_15919_ _13548_/A _13551_/X VGND VGND VPWR VPWR _15919_/Y sky130_fd_sc_hd__nor2_4
X_19687_ _19686_/Y _19682_/X _19612_/X _19682_/X VGND VGND VPWR VPWR _23664_/D sky130_fd_sc_hd__a2bb2o_4
X_16899_ _16147_/Y _24274_/Q _16147_/Y _24274_/Q VGND VGND VPWR VPWR _16899_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18638_ _18637_/Y VGND VGND VPWR VPWR _18805_/A sky130_fd_sc_hd__buf_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17972__B2 _17973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18569_ _18400_/Y _18568_/X VGND VGND VPWR VPWR _18569_/X sky130_fd_sc_hd__or2_4
XANTENNA__16195__A _16382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20600_ _14425_/A _18893_/A VGND VGND VPWR VPWR _20603_/B sky130_fd_sc_hd__or2_4
XFILLER_178_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21580_ _21580_/A VGND VGND VPWR VPWR _21580_/X sky130_fd_sc_hd__buf_2
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20531_ _20476_/D _20476_/B _20529_/X _20531_/D VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__or4_4
XFILLER_166_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22644__B _22789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23250_ _23250_/A _23183_/B VGND VGND VPWR VPWR _23253_/B sky130_fd_sc_hd__or2_4
X_20462_ _24099_/Q _20457_/X VGND VGND VPWR VPWR _20462_/X sky130_fd_sc_hd__and2_4
XFILLER_119_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15750__A3 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22201_ _22201_/A _21311_/A VGND VGND VPWR VPWR _22202_/B sky130_fd_sc_hd__or2_4
XFILLER_192_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23181_ _20808_/Y _23006_/X _20947_/Y _22808_/X VGND VGND VPWR VPWR _23181_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22481__B1 _22465_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20393_ _23408_/Q VGND VGND VPWR VPWR _21952_/B sky130_fd_sc_hd__inv_2
X_22132_ _14272_/Y _21375_/X _17432_/Y _21733_/B VGND VGND VPWR VPWR _22132_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16160__B1 _16066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22660__A _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22063_ _21386_/B VGND VGND VPWR VPWR _22524_/B sky130_fd_sc_hd__buf_2
XFILLER_245_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21014_ _21012_/Y _14804_/Y _21013_/C VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__or3_4
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23194__C _23187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17660__B1 _17611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22965_ _21427_/A _22963_/X _22844_/X _22964_/X VGND VGND VPWR VPWR _22966_/A sky130_fd_sc_hd__o22a_4
XFILLER_216_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24704_ _25444_/CLK _16131_/X HRESETn VGND VGND VPWR VPWR _22883_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21916_ _22228_/A _21916_/B _21915_/X VGND VGND VPWR VPWR _21916_/X sky130_fd_sc_hd__and3_4
XFILLER_55_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22896_ _16229_/A _23010_/B VGND VGND VPWR VPWR _22900_/B sky130_fd_sc_hd__or2_4
XFILLER_16_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14226__B1 _13809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21847_ _21847_/A VGND VGND VPWR VPWR _21847_/Y sky130_fd_sc_hd__inv_2
X_24635_ _24629_/CLK _16328_/X HRESETn VGND VGND VPWR VPWR _24635_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12579_/Y _24873_/Q _12579_/Y _24873_/Q VGND VGND VPWR VPWR _12587_/A sky130_fd_sc_hd__a2bb2o_4
X_24566_ _24566_/CLK _24566_/D HRESETn VGND VGND VPWR VPWR _16512_/A sky130_fd_sc_hd__dfrtp_4
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21778_ _21275_/A VGND VGND VPWR VPWR _22390_/A sky130_fd_sc_hd__buf_2
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _20728_/X VGND VGND VPWR VPWR _24022_/D sky130_fd_sc_hd__inv_2
X_23517_ _23918_/CLK _20098_/X VGND VGND VPWR VPWR _13453_/B sky130_fd_sc_hd__dfxtp_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24497_ _24532_/CLK _16698_/X HRESETn VGND VGND VPWR VPWR _16696_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_168_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _25199_/Q VGND VGND VPWR VPWR _14250_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23448_ _23529_/CLK _23448_/D VGND VGND VPWR VPWR _23448_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13197_/X _13200_/X _13183_/X VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__o21a_4
XFILLER_125_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14181_ _14181_/A VGND VGND VPWR VPWR _14181_/X sky130_fd_sc_hd__buf_2
X_23379_ _21022_/X VGND VGND VPWR VPWR IRQ[23] sky130_fd_sc_hd__buf_2
XANTENNA__18140__A1 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13132_ _13130_/Y _13132_/B VGND VGND VPWR VPWR _13132_/X sky130_fd_sc_hd__and2_4
X_25118_ _24095_/CLK _14508_/X HRESETn VGND VGND VPWR VPWR _25118_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16151__B1 _15905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13063_ _13068_/A _13063_/B _12312_/X _13066_/B VGND VGND VPWR VPWR _13069_/B sky130_fd_sc_hd__or4_4
X_17940_ _17944_/A _23884_/Q VGND VGND VPWR VPWR _17940_/X sky130_fd_sc_hd__or2_4
X_25049_ _24000_/CLK _14876_/X HRESETn VGND VGND VPWR VPWR _25049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12014_ _24105_/Q _12000_/X _12013_/Y VGND VGND VPWR VPWR _12015_/A sky130_fd_sc_hd__o21a_4
X_17871_ _17871_/A _17871_/B VGND VGND VPWR VPWR _17873_/B sky130_fd_sc_hd__or2_4
Xclkbuf_4_6_0_HCLK clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19610_ _19610_/A VGND VGND VPWR VPWR _19610_/X sky130_fd_sc_hd__buf_2
XFILLER_239_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16822_ _16822_/A VGND VGND VPWR VPWR _16822_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19541_ _19528_/Y VGND VGND VPWR VPWR _19541_/X sky130_fd_sc_hd__buf_2
X_16753_ _15051_/Y _16748_/X _16402_/X _16752_/X VGND VGND VPWR VPWR _24475_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13965_ _13934_/X VGND VGND VPWR VPWR _13967_/A sky130_fd_sc_hd__inv_2
XFILLER_207_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15704_ _15703_/X VGND VGND VPWR VPWR _15704_/X sky130_fd_sc_hd__buf_2
XFILLER_47_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22729__B _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12916_ _12857_/A _12915_/Y VGND VGND VPWR VPWR _12916_/X sky130_fd_sc_hd__or2_4
X_19472_ _18152_/B VGND VGND VPWR VPWR _19472_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16684_ _24502_/Q VGND VGND VPWR VPWR _16684_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14217__B1 _13806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _13896_/A VGND VGND VPWR VPWR _13924_/C sky130_fd_sc_hd__buf_2
XFILLER_62_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17004__A1_N _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18423_ _18423_/A VGND VGND VPWR VPWR _18476_/A sky130_fd_sc_hd__inv_2
X_15635_ _15626_/A VGND VGND VPWR VPWR _15635_/X sky130_fd_sc_hd__buf_2
XFILLER_206_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12847_ _12846_/X VGND VGND VPWR VPWR _12988_/A sky130_fd_sc_hd__buf_2
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18354_ _13199_/A _18347_/B _18351_/X VGND VGND VPWR VPWR _18354_/Y sky130_fd_sc_hd__a21oi_4
X_15566_ _15565_/X _15560_/X VGND VGND VPWR VPWR _15569_/A sky130_fd_sc_hd__or2_4
XFILLER_187_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16260__A1_N _16259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12778_ _24798_/Q VGND VGND VPWR VPWR _12778_/Y sky130_fd_sc_hd__inv_2
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15980__A3 _16245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18903__B1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17305_/A _17305_/B VGND VGND VPWR VPWR _17306_/C sky130_fd_sc_hd__or2_4
X_14517_ _14517_/A VGND VGND VPWR VPWR _14517_/Y sky130_fd_sc_hd__inv_2
X_11729_ _14199_/A _11728_/X VGND VGND VPWR VPWR _11729_/X sky130_fd_sc_hd__or2_4
X_18285_ _18283_/X _17713_/X _17723_/X _18285_/D VGND VGND VPWR VPWR _18285_/X sky130_fd_sc_hd__and4_4
X_15497_ _15496_/X VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__buf_2
XANTENNA__16743__A _16762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _24645_/Q _17227_/Y _16363_/Y _17250_/A VGND VGND VPWR VPWR _17236_/X sky130_fd_sc_hd__a2bb2o_4
X_14448_ _25141_/Q VGND VGND VPWR VPWR _14448_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23255__A2 _22673_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _17165_/Y _17167_/B _17160_/C VGND VGND VPWR VPWR _17167_/X sky130_fd_sc_hd__and3_4
XANTENNA__22463__B1 _16612_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24796__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14379_ _25160_/Q _14360_/A _25159_/Q _14354_/B VGND VGND VPWR VPWR _14379_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16118_ _23061_/A VGND VGND VPWR VPWR _16118_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16142__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24725__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17098_ _17097_/X VGND VGND VPWR VPWR _24400_/D sky130_fd_sc_hd__inv_2
Xclkbuf_8_151_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _24171_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17574__A _24312_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16049_ _16044_/A VGND VGND VPWR VPWR _16049_/X sky130_fd_sc_hd__buf_2
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17642__B1 _17611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19808_ _21621_/B _19806_/X _19807_/X _19806_/X VGND VGND VPWR VPWR _23623_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13607__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14456__B1 _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19739_ _19738_/Y _19733_/X _19620_/X _19719_/Y VGND VGND VPWR VPWR _23645_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19395__B1 _19305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22750_ _22750_/A VGND VGND VPWR VPWR _22750_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21701_ _23422_/Q _20344_/X _23398_/Q _21656_/X VGND VGND VPWR VPWR _21701_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22681_ _22681_/A VGND VGND VPWR VPWR _22681_/Y sky130_fd_sc_hd__inv_2
XFILLER_213_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24420_ _24425_/CLK _24420_/D HRESETn VGND VGND VPWR VPWR _24420_/Q sky130_fd_sc_hd__dfrtp_4
X_21632_ _14709_/X _21624_/X _21631_/X VGND VGND VPWR VPWR _21632_/X sky130_fd_sc_hd__or3_4
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12234__A2 _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24351_ _24625_/CLK _24351_/D HRESETn VGND VGND VPWR VPWR _24351_/Q sky130_fd_sc_hd__dfrtp_4
X_21563_ _21558_/X _21563_/B _21563_/C _21563_/D VGND VGND VPWR VPWR _21564_/B sky130_fd_sc_hd__and4_4
XANTENNA__17749__A _24293_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16653__A _16653_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23302_ _23302_/A _23301_/X _22150_/A VGND VGND VPWR VPWR _23302_/X sky130_fd_sc_hd__or3_4
XFILLER_178_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15484__A1_N _15482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20514_ _20470_/A _14073_/A _20463_/A _20514_/D VGND VGND VPWR VPWR _20514_/X sky130_fd_sc_hd__and4_4
X_24282_ _24283_/CLK _17830_/X HRESETn VGND VGND VPWR VPWR _24282_/Q sky130_fd_sc_hd__dfrtp_4
X_21494_ _21472_/A VGND VGND VPWR VPWR _21808_/A sky130_fd_sc_hd__buf_2
X_23233_ _23118_/X _23233_/B VGND VGND VPWR VPWR _23240_/C sky130_fd_sc_hd__and2_4
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11797__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20445_ _20445_/A _24099_/Q _24095_/Q VGND VGND VPWR VPWR _20445_/X sky130_fd_sc_hd__or3_4
XANTENNA__22454__B1 _25381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23164_ _23118_/X _23164_/B VGND VGND VPWR VPWR _23173_/C sky130_fd_sc_hd__and2_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16133__B1 _15972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20376_ _23414_/Q VGND VGND VPWR VPWR _21672_/B sky130_fd_sc_hd__inv_2
XANTENNA__22390__A _22390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22115_ _22115_/A VGND VGND VPWR VPWR _22115_/Y sky130_fd_sc_hd__inv_2
X_23095_ _12425_/A _23280_/A _23094_/X VGND VGND VPWR VPWR _23095_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22046_ _22032_/A _20328_/Y VGND VGND VPWR VPWR _22046_/X sky130_fd_sc_hd__or2_4
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14447__B1 _14420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ _23998_/CLK _23997_/D HRESETn VGND VGND VPWR VPWR _20668_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16828__A _16810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22549__B _22549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19386__B1 _19341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15732__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13750_ _24517_/Q _24516_/Q _24518_/Q VGND VGND VPWR VPWR _14775_/B sky130_fd_sc_hd__and3_4
X_22948_ _24470_/Q _22543_/A _22903_/X VGND VGND VPWR VPWR _22948_/X sky130_fd_sc_hd__o21a_4
XFILLER_216_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ _12730_/A VGND VGND VPWR VPWR _12728_/A sky130_fd_sc_hd__buf_2
X_13681_ _25304_/Q _13679_/X _13680_/Y VGND VGND VPWR VPWR _13681_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22879_ _22788_/X _22878_/X _22497_/X _24739_/Q _22498_/X VGND VGND VPWR VPWR _22880_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15420_ _15399_/X _15420_/B _15427_/C VGND VGND VPWR VPWR _24986_/D sky130_fd_sc_hd__and3_4
X_12632_ _12601_/Y _12702_/A _12631_/X VGND VGND VPWR VPWR _12633_/A sky130_fd_sc_hd__or3_4
X_24618_ _24485_/CLK _24618_/D HRESETn VGND VGND VPWR VPWR _24618_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _12563_/A VGND VGND VPWR VPWR _12619_/A sky130_fd_sc_hd__inv_2
X_15351_ _15347_/A _15346_/X VGND VGND VPWR VPWR _15351_/Y sky130_fd_sc_hd__nand2_4
XFILLER_157_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24549_ _24542_/CLK _24549_/D HRESETn VGND VGND VPWR VPWR _16558_/A sky130_fd_sc_hd__dfrtp_4
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14302_ _13531_/D _14301_/Y _14310_/A VGND VGND VPWR VPWR _25187_/D sky130_fd_sc_hd__o21a_4
X_18070_ _15704_/X _18050_/X _18069_/X _24253_/Q _18029_/X VGND VGND VPWR VPWR _18070_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_196_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12212_/X _12480_/X _12421_/A _12491_/B VGND VGND VPWR VPWR _12494_/X sky130_fd_sc_hd__a211o_4
X_15282_ _15282_/A _15282_/B VGND VGND VPWR VPWR _15283_/C sky130_fd_sc_hd__or2_4
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _16078_/Y _24381_/Q _24722_/Q _17053_/C VGND VGND VPWR VPWR _17021_/X sky130_fd_sc_hd__a2bb2o_4
X_14233_ _14233_/A VGND VGND VPWR VPWR _14233_/X sky130_fd_sc_hd__buf_2
XANTENNA__22445__B1 _11837_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19310__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14164_ _14155_/X _14163_/Y _25142_/Q _14155_/X VGND VGND VPWR VPWR _25222_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16124__B1 _15963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21909__A _22093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13115_ _13115_/A _13115_/B VGND VGND VPWR VPWR _13115_/X sky130_fd_sc_hd__or2_4
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_224_0_HCLK clkbuf_7_112_0_HCLK/X VGND VGND VPWR VPWR _25154_/CLK sky130_fd_sc_hd__clkbuf_1
X_14095_ _24013_/Q _14066_/A _14082_/X _14028_/A _14093_/X VGND VGND VPWR VPWR _25236_/D
+ sky130_fd_sc_hd__a32o_4
X_18972_ _18971_/Y _18966_/X _16796_/X _18966_/X VGND VGND VPWR VPWR _23912_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13046_ _12363_/A _13046_/B VGND VGND VPWR VPWR _13046_/X sky130_fd_sc_hd__or2_4
X_17923_ _15693_/A _14778_/X _15923_/X _17922_/X VGND VGND VPWR VPWR _17924_/B sky130_fd_sc_hd__a211o_4
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13427__A _13322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17854_ _17853_/X VGND VGND VPWR VPWR _17854_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14438__B1 _14248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16805_ _16857_/A VGND VGND VPWR VPWR _16805_/X sky130_fd_sc_hd__buf_2
XFILLER_208_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17785_ _16957_/X _17774_/X VGND VGND VPWR VPWR _17788_/B sky130_fd_sc_hd__or2_4
X_14997_ _14921_/X _16764_/A _14921_/X _16764_/A VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16738__A _16737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19524_ _23717_/Q VGND VGND VPWR VPWR _21199_/B sky130_fd_sc_hd__inv_2
XFILLER_35_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16736_ _24482_/Q VGND VGND VPWR VPWR _16736_/Y sky130_fd_sc_hd__inv_2
X_13948_ _13934_/X _13947_/Y _13948_/C _13899_/X VGND VGND VPWR VPWR _13949_/A sky130_fd_sc_hd__or4_4
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_223_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19455_ _19453_/Y _19451_/X _19454_/X _19451_/X VGND VGND VPWR VPWR _19455_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16667_ _16654_/X VGND VGND VPWR VPWR _16667_/X sky130_fd_sc_hd__buf_2
X_13879_ _13861_/X _13878_/X _14270_/A _13876_/X VGND VGND VPWR VPWR _25255_/D sky130_fd_sc_hd__o22a_4
XFILLER_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18406_ _22557_/A _18479_/D _16209_/Y _24189_/Q VGND VGND VPWR VPWR _18406_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15618_ _15618_/A VGND VGND VPWR VPWR _15618_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19386_ _19385_/Y _19382_/X _19341_/X _19382_/X VGND VGND VPWR VPWR _23766_/D sky130_fd_sc_hd__a2bb2o_4
X_16598_ _16596_/Y _16592_/X _16241_/X _16597_/X VGND VGND VPWR VPWR _24534_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22279__A3 _22274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18337_ _18334_/X _20079_/B _19119_/C VGND VGND VPWR VPWR _19815_/A sky130_fd_sc_hd__or3_4
X_15549_ _13603_/A VGND VGND VPWR VPWR _15549_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18268_ _18268_/A VGND VGND VPWR VPWR _18268_/X sky130_fd_sc_hd__buf_2
XFILLER_147_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24906__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17219_ _16338_/Y _24360_/Q _16338_/Y _24360_/Q VGND VGND VPWR VPWR _17219_/X sky130_fd_sc_hd__a2bb2o_4
X_18199_ _18199_/A _19205_/A VGND VGND VPWR VPWR _18201_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20230_ _23469_/Q VGND VGND VPWR VPWR _20230_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19852__B2 _19851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20161_ _21790_/B _20156_/X _20115_/X _20156_/X VGND VGND VPWR VPWR _23496_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12309__A2_N _24850_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20092_ _23519_/Q VGND VGND VPWR VPWR _20092_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23920_ _23918_/CLK _23920_/D VGND VGND VPWR VPWR _18949_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_84_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14429__B1 _14427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23851_ _23850_/CLK _23851_/D VGND VGND VPWR VPWR _23851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22802_ _22694_/B VGND VGND VPWR VPWR _22890_/B sky130_fd_sc_hd__buf_2
X_20994_ _20994_/A VGND VGND VPWR VPWR _20996_/A sky130_fd_sc_hd__inv_2
X_23782_ _24252_/CLK _19342_/X VGND VGND VPWR VPWR _18177_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_226_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25521_ _25520_/CLK _25521_/D HRESETn VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__dfrtp_4
X_22733_ _24767_/Q _22283_/X _15863_/X _24839_/Q _22444_/X VGND VGND VPWR VPWR _22733_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_213_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22664_ _23093_/A _22663_/X VGND VGND VPWR VPWR _22676_/B sky130_fd_sc_hd__and2_4
X_25452_ _25454_/CLK _12467_/Y HRESETn VGND VGND VPWR VPWR _12246_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15944__A3 HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21615_ _14766_/X VGND VGND VPWR VPWR _21648_/A sky130_fd_sc_hd__buf_2
X_24403_ _24952_/CLK _24403_/D HRESETn VGND VGND VPWR VPWR _24403_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_116_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22675__B1 _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22595_ _22595_/A _22595_/B VGND VGND VPWR VPWR _22595_/X sky130_fd_sc_hd__and2_4
X_25383_ _25402_/CLK _25383_/D HRESETn VGND VGND VPWR VPWR _25383_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16383__A _16390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21546_ _21545_/X VGND VGND VPWR VPWR _21546_/Y sky130_fd_sc_hd__inv_2
X_24334_ _24334_/CLK _24334_/D HRESETn VGND VGND VPWR VPWR _24334_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24647__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24265_ _24715_/CLK _17892_/X HRESETn VGND VGND VPWR VPWR _16929_/A sky130_fd_sc_hd__dfrtp_4
X_21477_ _21673_/A _21477_/B VGND VGND VPWR VPWR _21477_/X sky130_fd_sc_hd__or2_4
XFILLER_181_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23216_ _24042_/Q _21296_/X _24074_/Q _21320_/X VGND VGND VPWR VPWR _23216_/Y sky130_fd_sc_hd__a22oi_4
X_20428_ _20427_/Y _20423_/X _11851_/A _20423_/X VGND VGND VPWR VPWR _20428_/X sky130_fd_sc_hd__a2bb2o_4
X_24196_ _24196_/CLK _24196_/D HRESETn VGND VGND VPWR VPWR _24196_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16105__A1_N _16102_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23147_ _16212_/A _23183_/B VGND VGND VPWR VPWR _23147_/X sky130_fd_sc_hd__or2_4
X_20359_ _21991_/B _20352_/X _19832_/X _20352_/A VGND VGND VPWR VPWR _20359_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23078_ _16574_/A _22940_/X _22941_/X _23077_/X VGND VGND VPWR VPWR _23079_/C sky130_fd_sc_hd__a211o_4
XFILLER_103_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14920_ _14920_/A VGND VGND VPWR VPWR _14921_/A sky130_fd_sc_hd__inv_2
X_22029_ _22029_/A _22029_/B _22029_/C VGND VGND VPWR VPWR _22029_/X sky130_fd_sc_hd__and3_4
XANTENNA__17942__A _18023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_54_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24407_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ _14819_/X _14850_/X _25201_/Q _14844_/X VGND VGND VPWR VPWR _14851_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_248_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13802_ _13802_/A VGND VGND VPWR VPWR _21384_/B sky130_fd_sc_hd__buf_2
X_17570_ _24322_/Q VGND VGND VPWR VPWR _17610_/A sky130_fd_sc_hd__inv_2
X_14782_ _14781_/X VGND VGND VPWR VPWR _14785_/B sky130_fd_sc_hd__inv_2
XANTENNA__21166__B1 _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11994_ _11663_/A _11663_/B _11993_/Y VGND VGND VPWR VPWR _11994_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16521_ _16519_/Y _16520_/X _16252_/X _16520_/X VGND VGND VPWR VPWR _16521_/X sky130_fd_sc_hd__a2bb2o_4
X_13733_ _13695_/B _13732_/Y _13730_/X _13723_/X _11685_/A VGND VGND VPWR VPWR _25291_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_216_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19240_ _13274_/B VGND VGND VPWR VPWR _19240_/Y sky130_fd_sc_hd__inv_2
X_16452_ _15124_/Y _16446_/X _16451_/X _16446_/X VGND VGND VPWR VPWR _24587_/D sky130_fd_sc_hd__a2bb2o_4
X_13664_ _24050_/Q _13664_/B VGND VGND VPWR VPWR _13664_/X sky130_fd_sc_hd__or2_4
XANTENNA__16593__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22295__A _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15935__A3 _15933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15403_ _15120_/Y _15409_/B VGND VGND VPWR VPWR _15407_/B sky130_fd_sc_hd__or2_4
X_12615_ _25434_/Q VGND VGND VPWR VPWR _12642_/A sky130_fd_sc_hd__inv_2
X_19171_ _23843_/Q VGND VGND VPWR VPWR _19171_/Y sky130_fd_sc_hd__inv_2
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22726__C _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17389__A _17389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16383_ _16390_/A VGND VGND VPWR VPWR _16384_/A sky130_fd_sc_hd__buf_2
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22666__B1 _24838_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13595_ _13857_/A _14569_/B _13840_/A _14601_/A VGND VGND VPWR VPWR _13595_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18122_ _17975_/X _18120_/X _18122_/C VGND VGND VPWR VPWR _18123_/C sky130_fd_sc_hd__and3_4
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15334_ _15096_/Y _15316_/X _15340_/A _15334_/D VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__or4_4
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12546_ _25414_/Q _12545_/A _12725_/A _12545_/Y VGND VGND VPWR VPWR _12553_/B sky130_fd_sc_hd__o22a_4
X_18053_ _18126_/A _19060_/A VGND VGND VPWR VPWR _18054_/C sky130_fd_sc_hd__or2_4
XFILLER_177_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15265_ _15271_/A _15268_/A _15259_/X VGND VGND VPWR VPWR _15265_/X sky130_fd_sc_hd__or3_4
X_12477_ _12205_/Y _12391_/X VGND VGND VPWR VPWR _12478_/B sky130_fd_sc_hd__or2_4
XFILLER_138_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17004_ _24722_/Q _17053_/C _24726_/Q _17139_/A VGND VGND VPWR VPWR _17004_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14216_ _20497_/B VGND VGND VPWR VPWR _20525_/B sky130_fd_sc_hd__inv_2
XANTENNA__21639__A _22388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15196_ _15196_/A _15193_/X VGND VGND VPWR VPWR _15197_/C sky130_fd_sc_hd__or2_4
XFILLER_153_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ _14134_/X _14146_/Y _14112_/A _14134_/X VGND VGND VPWR VPWR _14147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_193_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18013__A _18013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14078_ _14066_/A VGND VGND VPWR VPWR _14078_/X sky130_fd_sc_hd__buf_2
X_18955_ _18954_/Y _18952_/X _18908_/X _18952_/X VGND VGND VPWR VPWR _23918_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22197__A2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13029_ _13021_/C _13021_/D VGND VGND VPWR VPWR _13029_/X sky130_fd_sc_hd__or2_4
X_17906_ _17903_/Y _17913_/B _17905_/Y VGND VGND VPWR VPWR _17907_/B sky130_fd_sc_hd__o21ai_4
XFILLER_239_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18886_ _23959_/Q _18886_/B VGND VGND VPWR VPWR _18887_/B sky130_fd_sc_hd__or2_4
XANTENNA__23952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ _17852_/A _17832_/X _17836_/X VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__and3_4
XFILLER_55_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16468__A _16468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17768_ _16914_/Y _17832_/A _16923_/Y _17768_/D VGND VGND VPWR VPWR _17769_/D sky130_fd_sc_hd__or4_4
XFILLER_208_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16719_ _16718_/Y _16716_/X _16364_/X _16716_/X VGND VGND VPWR VPWR _24488_/D sky130_fd_sc_hd__a2bb2o_4
X_19507_ _19507_/A VGND VGND VPWR VPWR _19507_/Y sky130_fd_sc_hd__inv_2
X_17699_ _17529_/Y _17703_/B VGND VGND VPWR VPWR _17701_/B sky130_fd_sc_hd__or2_4
XANTENNA__19770__B1 _19769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19438_ _19438_/A VGND VGND VPWR VPWR _19438_/X sky130_fd_sc_hd__buf_2
XFILLER_211_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19369_ _19368_/Y VGND VGND VPWR VPWR _19369_/X sky130_fd_sc_hd__buf_2
XFILLER_10_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21400_ _21408_/A _21400_/B VGND VGND VPWR VPWR _21401_/C sky130_fd_sc_hd__or2_4
XFILLER_210_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13620__A _18098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22380_ _22380_/A _22380_/B _22379_/X VGND VGND VPWR VPWR _22380_/X sky130_fd_sc_hd__and3_4
XANTENNA__24740__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22933__A _16003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21331_ _21574_/A VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__buf_2
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24050_ _24488_/CLK _20849_/Y HRESETn VGND VGND VPWR VPWR _24050_/Q sky130_fd_sc_hd__dfrtp_4
X_21262_ _21262_/A _21252_/X _21261_/X VGND VGND VPWR VPWR _21262_/X sky130_fd_sc_hd__or3_4
XANTENNA__21549__A _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23001_ _22999_/X _23000_/X _22929_/X VGND VGND VPWR VPWR _23001_/X sky130_fd_sc_hd__or3_4
X_20213_ _20213_/A VGND VGND VPWR VPWR _20213_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15547__A _15544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21193_ _21204_/A _21190_/X _21193_/C VGND VGND VPWR VPWR _21193_/X sky130_fd_sc_hd__and3_4
XFILLER_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20144_ _21403_/B _20141_/X _20122_/X _20141_/X VGND VGND VPWR VPWR _23502_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20075_ _20074_/Y _20072_/X _19810_/X _20072_/X VGND VGND VPWR VPWR _23526_/D sky130_fd_sc_hd__a2bb2o_4
X_24952_ _24952_/CLK _15504_/X HRESETn VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__20199__B2 _20198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23903_ _25082_/CLK _23903_/D VGND VGND VPWR VPWR _18994_/A sky130_fd_sc_hd__dfxtp_4
X_24883_ _24883_/CLK _24883_/D HRESETn VGND VGND VPWR VPWR _24883_/Q sky130_fd_sc_hd__dfrtp_4
X_23834_ _23830_/CLK _19197_/X VGND VGND VPWR VPWR _19195_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_245_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13086__C1 _13040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19689__A _19675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20977_ _20977_/A _13529_/A VGND VGND VPWR VPWR _20977_/X sky130_fd_sc_hd__and2_4
X_23765_ _23768_/CLK _23765_/D VGND VGND VPWR VPWR _18206_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24899__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25504_ _25507_/CLK _11989_/X HRESETn VGND VGND VPWR VPWR _11662_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_26_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22716_ _22716_/A _22316_/B VGND VGND VPWR VPWR _22719_/B sky130_fd_sc_hd__or2_4
XANTENNA__24828__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16575__B1 _16315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23696_ _23407_/CLK _23696_/D VGND VGND VPWR VPWR _23696_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25435_ _25419_/CLK _12646_/X HRESETn VGND VGND VPWR VPWR _12644_/A sky130_fd_sc_hd__dfrtp_4
X_22647_ _22289_/A _22646_/X _21314_/X _16053_/A _21317_/X VGND VGND VPWR VPWR _22647_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_213_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12400_ _12393_/A _12400_/B VGND VGND VPWR VPWR _12401_/C sky130_fd_sc_hd__or2_4
X_13380_ _13412_/A _13378_/X _13379_/X VGND VGND VPWR VPWR _13384_/B sky130_fd_sc_hd__and3_4
XANTENNA__24481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22578_ _16703_/Y _22578_/B VGND VGND VPWR VPWR _22578_/X sky130_fd_sc_hd__and2_4
X_25366_ _25365_/CLK _25366_/D HRESETn VGND VGND VPWR VPWR _25366_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20123__B2 _20118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22663__A3 _22148_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12331_ _12329_/A _24849_/Q _12329_/Y _12330_/Y VGND VGND VPWR VPWR _12335_/C sky130_fd_sc_hd__o22a_4
X_24317_ _25543_/CLK _24317_/D HRESETn VGND VGND VPWR VPWR _17511_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16878__B2 _16877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21871__A1 _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21529_ _21231_/A VGND VGND VPWR VPWR _22721_/B sky130_fd_sc_hd__buf_2
XFILLER_127_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25297_ _25292_/CLK _25297_/D HRESETn VGND VGND VPWR VPWR _11666_/A sky130_fd_sc_hd__dfrtp_4
X_12262_ _12261_/Y _24775_/Q _25448_/Q _12199_/Y VGND VGND VPWR VPWR _12262_/X sky130_fd_sc_hd__a2bb2o_4
X_15050_ _25019_/Q _15037_/Y _14895_/X _24462_/Q VGND VGND VPWR VPWR _15056_/A sky130_fd_sc_hd__a2bb2o_4
X_24248_ _23754_/CLK _24248_/D HRESETn VGND VGND VPWR VPWR _24248_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16674__A1_N _16671_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15550__B2 _15547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14001_ _25244_/Q _13998_/X _14021_/D VGND VGND VPWR VPWR _14001_/X sky130_fd_sc_hd__or3_4
XANTENNA__12364__B2 _24848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12193_ _25463_/Q VGND VGND VPWR VPWR _12428_/A sky130_fd_sc_hd__inv_2
X_24179_ _24523_/CLK _24179_/D HRESETn VGND VGND VPWR VPWR _24179_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18740_ _18714_/A VGND VGND VPWR VPWR _18740_/X sky130_fd_sc_hd__buf_2
XFILLER_163_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15853__A2 _15774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15952_ HWDATA[27] VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__buf_2
XFILLER_209_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14903_ _14902_/Y VGND VGND VPWR VPWR _15206_/A sky130_fd_sc_hd__buf_2
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18671_ _16562_/A _18717_/A _16622_/Y _24135_/Q VGND VGND VPWR VPWR _18673_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15883_ _15858_/X _15865_/X _15734_/X _23119_/A _15872_/X VGND VGND VPWR VPWR _24815_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_209_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16288__A _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17622_ _17571_/Y _17621_/X VGND VGND VPWR VPWR _17626_/B sky130_fd_sc_hd__or2_4
X_14834_ _14852_/A VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__buf_2
XANTENNA__16802__B2 _16738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17553_ _17553_/A VGND VGND VPWR VPWR _17553_/Y sky130_fd_sc_hd__inv_2
X_14765_ _21248_/A VGND VGND VPWR VPWR _14765_/X sky130_fd_sc_hd__buf_2
X_11977_ _11713_/A _11968_/X _11975_/Y _25506_/Q _11976_/X VGND VGND VPWR VPWR _11977_/X
+ sky130_fd_sc_hd__o32a_4
X_16504_ _24569_/Q VGND VGND VPWR VPWR _16504_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13716_ _13688_/Y VGND VGND VPWR VPWR _13716_/X sky130_fd_sc_hd__buf_2
XFILLER_205_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17484_ _17484_/A _18333_/B _17484_/C _17484_/D VGND VGND VPWR VPWR _17484_/X sky130_fd_sc_hd__or4_4
XANTENNA__24569__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _21240_/A VGND VGND VPWR VPWR _21263_/A sky130_fd_sc_hd__buf_2
X_19223_ _19222_/Y _19217_/X _19131_/X _19217_/X VGND VGND VPWR VPWR _23824_/D sky130_fd_sc_hd__a2bb2o_4
X_16435_ _16442_/A VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__buf_2
XFILLER_176_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13647_ _13647_/A VGND VGND VPWR VPWR _13647_/X sky130_fd_sc_hd__buf_2
XANTENNA__22103__A2 _21091_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18008__A _18008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23300__B2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19154_ _23849_/Q VGND VGND VPWR VPWR _19154_/Y sky130_fd_sc_hd__inv_2
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16366_ _16363_/Y _16359_/X _16364_/X _16365_/X VGND VGND VPWR VPWR _24621_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16318__B1 _15960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13578_ _13578_/A VGND VGND VPWR VPWR _13578_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18105_ _18169_/A _18103_/X _18104_/X VGND VGND VPWR VPWR _18105_/X sky130_fd_sc_hd__and3_4
XFILLER_185_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15317_ _15096_/Y _15316_/X VGND VGND VPWR VPWR _15337_/B sky130_fd_sc_hd__or2_4
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _25422_/Q VGND VGND VPWR VPWR _12529_/Y sky130_fd_sc_hd__inv_2
X_19085_ _19085_/A VGND VGND VPWR VPWR _19085_/X sky130_fd_sc_hd__buf_2
X_16297_ _16290_/A VGND VGND VPWR VPWR _16325_/A sky130_fd_sc_hd__buf_2
XANTENNA__12056__A _14199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18036_ _18036_/A _23762_/Q VGND VGND VPWR VPWR _18036_/X sky130_fd_sc_hd__or2_4
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15248_ _15248_/A _15247_/X VGND VGND VPWR VPWR _15249_/A sky130_fd_sc_hd__or2_4
XANTENNA__15541__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15179_ _15068_/X _15177_/X _15178_/X VGND VGND VPWR VPWR _25044_/D sky130_fd_sc_hd__and3_4
XFILLER_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19987_ _17717_/X _18293_/X _19527_/C _19986_/X VGND VGND VPWR VPWR _19988_/A sky130_fd_sc_hd__or4_4
XFILLER_113_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _18938_/A _18938_/B _18938_/C VGND VGND VPWR VPWR _18938_/X sky130_fd_sc_hd__or3_4
.ends

