magic
tech sky130A
magscale 1 2
timestamp 1609941244
<< obsli1 >>
rect 1104 2159 118864 157777
<< obsm1 >>
rect 566 2128 119310 157808
<< metal2 >>
rect 1674 159200 1730 160000
rect 4802 159200 4858 160000
rect 7930 159200 7986 160000
rect 11058 159200 11114 160000
rect 14186 159200 14242 160000
rect 17130 159200 17186 160000
rect 20258 159200 20314 160000
rect 23386 159200 23442 160000
rect 26514 159200 26570 160000
rect 29642 159200 29698 160000
rect 32586 159200 32642 160000
rect 35714 159200 35770 160000
rect 38842 159200 38898 160000
rect 41970 159200 42026 160000
rect 45098 159200 45154 160000
rect 48226 159200 48282 160000
rect 51170 159200 51226 160000
rect 54298 159200 54354 160000
rect 57426 159200 57482 160000
rect 60554 159200 60610 160000
rect 63682 159200 63738 160000
rect 66810 159200 66866 160000
rect 69754 159200 69810 160000
rect 72882 159200 72938 160000
rect 76010 159200 76066 160000
rect 79138 159200 79194 160000
rect 82266 159200 82322 160000
rect 85210 159200 85266 160000
rect 88338 159200 88394 160000
rect 91466 159200 91522 160000
rect 94594 159200 94650 160000
rect 97722 159200 97778 160000
rect 100850 159200 100906 160000
rect 103794 159200 103850 160000
rect 106922 159200 106978 160000
rect 110050 159200 110106 160000
rect 113178 159200 113234 160000
rect 116306 159200 116362 160000
rect 119250 159200 119306 160000
rect 570 0 626 800
rect 3514 0 3570 800
rect 6642 0 6698 800
rect 9770 0 9826 800
rect 12898 0 12954 800
rect 16026 0 16082 800
rect 18970 0 19026 800
rect 22098 0 22154 800
rect 25226 0 25282 800
rect 28354 0 28410 800
rect 31482 0 31538 800
rect 34610 0 34666 800
rect 37554 0 37610 800
rect 40682 0 40738 800
rect 43810 0 43866 800
rect 46938 0 46994 800
rect 50066 0 50122 800
rect 53010 0 53066 800
rect 56138 0 56194 800
rect 59266 0 59322 800
rect 62394 0 62450 800
rect 65522 0 65578 800
rect 68650 0 68706 800
rect 71594 0 71650 800
rect 74722 0 74778 800
rect 77850 0 77906 800
rect 80978 0 81034 800
rect 84106 0 84162 800
rect 87234 0 87290 800
rect 90178 0 90234 800
rect 93306 0 93362 800
rect 96434 0 96490 800
rect 99562 0 99618 800
rect 102690 0 102746 800
rect 105634 0 105690 800
rect 108762 0 108818 800
rect 111890 0 111946 800
rect 115018 0 115074 800
rect 118146 0 118202 800
<< obsm2 >>
rect 572 159144 1618 159202
rect 1786 159144 4746 159202
rect 4914 159144 7874 159202
rect 8042 159144 11002 159202
rect 11170 159144 14130 159202
rect 14298 159144 17074 159202
rect 17242 159144 20202 159202
rect 20370 159144 23330 159202
rect 23498 159144 26458 159202
rect 26626 159144 29586 159202
rect 29754 159144 32530 159202
rect 32698 159144 35658 159202
rect 35826 159144 38786 159202
rect 38954 159144 41914 159202
rect 42082 159144 45042 159202
rect 45210 159144 48170 159202
rect 48338 159144 51114 159202
rect 51282 159144 54242 159202
rect 54410 159144 57370 159202
rect 57538 159144 60498 159202
rect 60666 159144 63626 159202
rect 63794 159144 66754 159202
rect 66922 159144 69698 159202
rect 69866 159144 72826 159202
rect 72994 159144 75954 159202
rect 76122 159144 79082 159202
rect 79250 159144 82210 159202
rect 82378 159144 85154 159202
rect 85322 159144 88282 159202
rect 88450 159144 91410 159202
rect 91578 159144 94538 159202
rect 94706 159144 97666 159202
rect 97834 159144 100794 159202
rect 100962 159144 103738 159202
rect 103906 159144 106866 159202
rect 107034 159144 109994 159202
rect 110162 159144 113122 159202
rect 113290 159144 116250 159202
rect 116418 159144 119194 159202
rect 572 856 119304 159144
rect 682 800 3458 856
rect 3626 800 6586 856
rect 6754 800 9714 856
rect 9882 800 12842 856
rect 13010 800 15970 856
rect 16138 800 18914 856
rect 19082 800 22042 856
rect 22210 800 25170 856
rect 25338 800 28298 856
rect 28466 800 31426 856
rect 31594 800 34554 856
rect 34722 800 37498 856
rect 37666 800 40626 856
rect 40794 800 43754 856
rect 43922 800 46882 856
rect 47050 800 50010 856
rect 50178 800 52954 856
rect 53122 800 56082 856
rect 56250 800 59210 856
rect 59378 800 62338 856
rect 62506 800 65466 856
rect 65634 800 68594 856
rect 68762 800 71538 856
rect 71706 800 74666 856
rect 74834 800 77794 856
rect 77962 800 80922 856
rect 81090 800 84050 856
rect 84218 800 87178 856
rect 87346 800 90122 856
rect 90290 800 93250 856
rect 93418 800 96378 856
rect 96546 800 99506 856
rect 99674 800 102634 856
rect 102802 800 105578 856
rect 105746 800 108706 856
rect 108874 800 111834 856
rect 112002 800 114962 856
rect 115130 800 118090 856
rect 118258 800 119304 856
<< metal3 >>
rect 0 156136 800 156256
rect 119200 154504 120000 154624
rect 0 151784 800 151904
rect 119200 149880 120000 150000
rect 0 147160 800 147280
rect 119200 145256 120000 145376
rect 0 142536 800 142656
rect 119200 140632 120000 140752
rect 0 137912 800 138032
rect 119200 136008 120000 136128
rect 0 133288 800 133408
rect 119200 131656 120000 131776
rect 0 128936 800 129056
rect 119200 127032 120000 127152
rect 0 124312 800 124432
rect 119200 122408 120000 122528
rect 0 119688 800 119808
rect 119200 117784 120000 117904
rect 0 115064 800 115184
rect 119200 113160 120000 113280
rect 0 110440 800 110560
rect 119200 108536 120000 108656
rect 0 105816 800 105936
rect 119200 104184 120000 104304
rect 0 101464 800 101584
rect 119200 99560 120000 99680
rect 0 96840 800 96960
rect 119200 94936 120000 95056
rect 0 92216 800 92336
rect 119200 90312 120000 90432
rect 0 87592 800 87712
rect 119200 85688 120000 85808
rect 0 82968 800 83088
rect 119200 81336 120000 81456
rect 0 78344 800 78464
rect 119200 76712 120000 76832
rect 0 73992 800 74112
rect 119200 72088 120000 72208
rect 0 69368 800 69488
rect 119200 67464 120000 67584
rect 0 64744 800 64864
rect 119200 62840 120000 62960
rect 0 60120 800 60240
rect 119200 58216 120000 58336
rect 0 55496 800 55616
rect 119200 53864 120000 53984
rect 0 51144 800 51264
rect 119200 49240 120000 49360
rect 0 46520 800 46640
rect 119200 44616 120000 44736
rect 0 41896 800 42016
rect 119200 39992 120000 40112
rect 0 37272 800 37392
rect 119200 35368 120000 35488
rect 0 32648 800 32768
rect 119200 30744 120000 30864
rect 0 28024 800 28144
rect 119200 26392 120000 26512
rect 0 23672 800 23792
rect 119200 21768 120000 21888
rect 0 19048 800 19168
rect 119200 17144 120000 17264
rect 0 14424 800 14544
rect 119200 12520 120000 12640
rect 0 9800 800 9920
rect 119200 7896 120000 8016
rect 0 5176 800 5296
rect 119200 3544 120000 3664
<< obsm3 >>
rect 798 156336 119200 157793
rect 880 156056 119200 156336
rect 798 154704 119200 156056
rect 798 154424 119120 154704
rect 798 151984 119200 154424
rect 880 151704 119200 151984
rect 798 150080 119200 151704
rect 798 149800 119120 150080
rect 798 147360 119200 149800
rect 880 147080 119200 147360
rect 798 145456 119200 147080
rect 798 145176 119120 145456
rect 798 142736 119200 145176
rect 880 142456 119200 142736
rect 798 140832 119200 142456
rect 798 140552 119120 140832
rect 798 138112 119200 140552
rect 880 137832 119200 138112
rect 798 136208 119200 137832
rect 798 135928 119120 136208
rect 798 133488 119200 135928
rect 880 133208 119200 133488
rect 798 131856 119200 133208
rect 798 131576 119120 131856
rect 798 129136 119200 131576
rect 880 128856 119200 129136
rect 798 127232 119200 128856
rect 798 126952 119120 127232
rect 798 124512 119200 126952
rect 880 124232 119200 124512
rect 798 122608 119200 124232
rect 798 122328 119120 122608
rect 798 119888 119200 122328
rect 880 119608 119200 119888
rect 798 117984 119200 119608
rect 798 117704 119120 117984
rect 798 115264 119200 117704
rect 880 114984 119200 115264
rect 798 113360 119200 114984
rect 798 113080 119120 113360
rect 798 110640 119200 113080
rect 880 110360 119200 110640
rect 798 108736 119200 110360
rect 798 108456 119120 108736
rect 798 106016 119200 108456
rect 880 105736 119200 106016
rect 798 104384 119200 105736
rect 798 104104 119120 104384
rect 798 101664 119200 104104
rect 880 101384 119200 101664
rect 798 99760 119200 101384
rect 798 99480 119120 99760
rect 798 97040 119200 99480
rect 880 96760 119200 97040
rect 798 95136 119200 96760
rect 798 94856 119120 95136
rect 798 92416 119200 94856
rect 880 92136 119200 92416
rect 798 90512 119200 92136
rect 798 90232 119120 90512
rect 798 87792 119200 90232
rect 880 87512 119200 87792
rect 798 85888 119200 87512
rect 798 85608 119120 85888
rect 798 83168 119200 85608
rect 880 82888 119200 83168
rect 798 81536 119200 82888
rect 798 81256 119120 81536
rect 798 78544 119200 81256
rect 880 78264 119200 78544
rect 798 76912 119200 78264
rect 798 76632 119120 76912
rect 798 74192 119200 76632
rect 880 73912 119200 74192
rect 798 72288 119200 73912
rect 798 72008 119120 72288
rect 798 69568 119200 72008
rect 880 69288 119200 69568
rect 798 67664 119200 69288
rect 798 67384 119120 67664
rect 798 64944 119200 67384
rect 880 64664 119200 64944
rect 798 63040 119200 64664
rect 798 62760 119120 63040
rect 798 60320 119200 62760
rect 880 60040 119200 60320
rect 798 58416 119200 60040
rect 798 58136 119120 58416
rect 798 55696 119200 58136
rect 880 55416 119200 55696
rect 798 54064 119200 55416
rect 798 53784 119120 54064
rect 798 51344 119200 53784
rect 880 51064 119200 51344
rect 798 49440 119200 51064
rect 798 49160 119120 49440
rect 798 46720 119200 49160
rect 880 46440 119200 46720
rect 798 44816 119200 46440
rect 798 44536 119120 44816
rect 798 42096 119200 44536
rect 880 41816 119200 42096
rect 798 40192 119200 41816
rect 798 39912 119120 40192
rect 798 37472 119200 39912
rect 880 37192 119200 37472
rect 798 35568 119200 37192
rect 798 35288 119120 35568
rect 798 32848 119200 35288
rect 880 32568 119200 32848
rect 798 30944 119200 32568
rect 798 30664 119120 30944
rect 798 28224 119200 30664
rect 880 27944 119200 28224
rect 798 26592 119200 27944
rect 798 26312 119120 26592
rect 798 23872 119200 26312
rect 880 23592 119200 23872
rect 798 21968 119200 23592
rect 798 21688 119120 21968
rect 798 19248 119200 21688
rect 880 18968 119200 19248
rect 798 17344 119200 18968
rect 798 17064 119120 17344
rect 798 14624 119200 17064
rect 880 14344 119200 14624
rect 798 12720 119200 14344
rect 798 12440 119120 12720
rect 798 10000 119200 12440
rect 880 9720 119200 10000
rect 798 8096 119200 9720
rect 798 7816 119120 8096
rect 798 5376 119200 7816
rect 880 5096 119200 5376
rect 798 3744 119200 5096
rect 798 3464 119120 3744
rect 798 851 119200 3464
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< obsm4 >>
rect 2635 2483 4128 157453
rect 4608 2483 19488 157453
rect 19968 2483 34848 157453
rect 35328 2483 50208 157453
rect 50688 2483 65568 157453
rect 66048 2483 80928 157453
rect 81408 2483 96288 157453
rect 96768 2483 111648 157453
rect 112128 2483 117333 157453
<< labels >>
rlabel metal3 s 119200 49240 120000 49360 6 EXT_IRQ
port 1 nsew signal input
rlabel metal2 s 29642 159200 29698 160000 6 HADDR[0]
port 2 nsew signal output
rlabel metal2 s 116306 159200 116362 160000 6 HADDR[10]
port 3 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 HADDR[11]
port 4 nsew signal output
rlabel metal2 s 54298 159200 54354 160000 6 HADDR[12]
port 5 nsew signal output
rlabel metal2 s 4802 159200 4858 160000 6 HADDR[13]
port 6 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 HADDR[14]
port 7 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 HADDR[15]
port 8 nsew signal output
rlabel metal3 s 119200 44616 120000 44736 6 HADDR[16]
port 9 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 HADDR[17]
port 10 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 HADDR[18]
port 11 nsew signal output
rlabel metal3 s 119200 21768 120000 21888 6 HADDR[19]
port 12 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 HADDR[1]
port 13 nsew signal output
rlabel metal3 s 119200 72088 120000 72208 6 HADDR[20]
port 14 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 HADDR[21]
port 15 nsew signal output
rlabel metal2 s 85210 159200 85266 160000 6 HADDR[22]
port 16 nsew signal output
rlabel metal2 s 119250 159200 119306 160000 6 HADDR[23]
port 17 nsew signal output
rlabel metal3 s 119200 39992 120000 40112 6 HADDR[24]
port 18 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 HADDR[25]
port 19 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 HADDR[26]
port 20 nsew signal output
rlabel metal3 s 119200 140632 120000 140752 6 HADDR[27]
port 21 nsew signal output
rlabel metal3 s 119200 3544 120000 3664 6 HADDR[28]
port 22 nsew signal output
rlabel metal3 s 119200 67464 120000 67584 6 HADDR[29]
port 23 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 HADDR[2]
port 24 nsew signal output
rlabel metal2 s 20258 159200 20314 160000 6 HADDR[30]
port 25 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 HADDR[31]
port 26 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 HADDR[3]
port 27 nsew signal output
rlabel metal3 s 119200 104184 120000 104304 6 HADDR[4]
port 28 nsew signal output
rlabel metal2 s 91466 159200 91522 160000 6 HADDR[5]
port 29 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 HADDR[6]
port 30 nsew signal output
rlabel metal3 s 119200 90312 120000 90432 6 HADDR[7]
port 31 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 HADDR[8]
port 32 nsew signal output
rlabel metal3 s 119200 127032 120000 127152 6 HADDR[9]
port 33 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 HCLK
port 34 nsew signal input
rlabel metal3 s 119200 108536 120000 108656 6 HRDATA[0]
port 35 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 HRDATA[10]
port 36 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 HRDATA[11]
port 37 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 HRDATA[12]
port 38 nsew signal input
rlabel metal2 s 26514 159200 26570 160000 6 HRDATA[13]
port 39 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 HRDATA[14]
port 40 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 HRDATA[15]
port 41 nsew signal input
rlabel metal3 s 119200 35368 120000 35488 6 HRDATA[16]
port 42 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 HRDATA[17]
port 43 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 HRDATA[18]
port 44 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 HRDATA[19]
port 45 nsew signal input
rlabel metal3 s 119200 53864 120000 53984 6 HRDATA[1]
port 46 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 HRDATA[20]
port 47 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 HRDATA[21]
port 48 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 HRDATA[22]
port 49 nsew signal input
rlabel metal2 s 100850 159200 100906 160000 6 HRDATA[23]
port 50 nsew signal input
rlabel metal3 s 119200 81336 120000 81456 6 HRDATA[24]
port 51 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 HRDATA[25]
port 52 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 HRDATA[26]
port 53 nsew signal input
rlabel metal3 s 119200 58216 120000 58336 6 HRDATA[27]
port 54 nsew signal input
rlabel metal3 s 119200 12520 120000 12640 6 HRDATA[28]
port 55 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 HRDATA[29]
port 56 nsew signal input
rlabel metal2 s 14186 159200 14242 160000 6 HRDATA[2]
port 57 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 HRDATA[30]
port 58 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 HRDATA[31]
port 59 nsew signal input
rlabel metal3 s 119200 113160 120000 113280 6 HRDATA[3]
port 60 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 HRDATA[4]
port 61 nsew signal input
rlabel metal2 s 17130 159200 17186 160000 6 HRDATA[5]
port 62 nsew signal input
rlabel metal2 s 45098 159200 45154 160000 6 HRDATA[6]
port 63 nsew signal input
rlabel metal2 s 1674 159200 1730 160000 6 HRDATA[7]
port 64 nsew signal input
rlabel metal3 s 119200 149880 120000 150000 6 HRDATA[8]
port 65 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 HRDATA[9]
port 66 nsew signal input
rlabel metal2 s 51170 159200 51226 160000 6 HREADY
port 67 nsew signal input
rlabel metal3 s 119200 62840 120000 62960 6 HRESETn
port 68 nsew signal input
rlabel metal2 s 72882 159200 72938 160000 6 HSIZE[0]
port 69 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 HSIZE[1]
port 70 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 HSIZE[2]
port 71 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 HTRANS[0]
port 72 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 HTRANS[1]
port 73 nsew signal output
rlabel metal2 s 82266 159200 82322 160000 6 HWDATA[0]
port 74 nsew signal output
rlabel metal2 s 63682 159200 63738 160000 6 HWDATA[10]
port 75 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 HWDATA[11]
port 76 nsew signal output
rlabel metal3 s 119200 85688 120000 85808 6 HWDATA[12]
port 77 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 HWDATA[13]
port 78 nsew signal output
rlabel metal3 s 119200 26392 120000 26512 6 HWDATA[14]
port 79 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 HWDATA[15]
port 80 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 HWDATA[16]
port 81 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 HWDATA[17]
port 82 nsew signal output
rlabel metal2 s 11058 159200 11114 160000 6 HWDATA[18]
port 83 nsew signal output
rlabel metal2 s 76010 159200 76066 160000 6 HWDATA[19]
port 84 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 HWDATA[1]
port 85 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 HWDATA[20]
port 86 nsew signal output
rlabel metal3 s 119200 136008 120000 136128 6 HWDATA[21]
port 87 nsew signal output
rlabel metal3 s 119200 7896 120000 8016 6 HWDATA[22]
port 88 nsew signal output
rlabel metal2 s 35714 159200 35770 160000 6 HWDATA[23]
port 89 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 HWDATA[24]
port 90 nsew signal output
rlabel metal3 s 119200 17144 120000 17264 6 HWDATA[25]
port 91 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 HWDATA[26]
port 92 nsew signal output
rlabel metal2 s 66810 159200 66866 160000 6 HWDATA[27]
port 93 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 HWDATA[28]
port 94 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 HWDATA[29]
port 95 nsew signal output
rlabel metal3 s 119200 131656 120000 131776 6 HWDATA[2]
port 96 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 HWDATA[30]
port 97 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 HWDATA[31]
port 98 nsew signal output
rlabel metal2 s 69754 159200 69810 160000 6 HWDATA[3]
port 99 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 HWDATA[4]
port 100 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 HWDATA[5]
port 101 nsew signal output
rlabel metal2 s 97722 159200 97778 160000 6 HWDATA[6]
port 102 nsew signal output
rlabel metal2 s 88338 159200 88394 160000 6 HWDATA[7]
port 103 nsew signal output
rlabel metal2 s 94594 159200 94650 160000 6 HWDATA[8]
port 104 nsew signal output
rlabel metal3 s 0 151784 800 151904 6 HWDATA[9]
port 105 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 HWRITE
port 106 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 IRQ[0]
port 107 nsew signal input
rlabel metal2 s 570 0 626 800 6 IRQ[10]
port 108 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 IRQ[11]
port 109 nsew signal input
rlabel metal2 s 7930 159200 7986 160000 6 IRQ[12]
port 110 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 IRQ[13]
port 111 nsew signal input
rlabel metal3 s 119200 30744 120000 30864 6 IRQ[14]
port 112 nsew signal input
rlabel metal2 s 38842 159200 38898 160000 6 IRQ[1]
port 113 nsew signal input
rlabel metal2 s 48226 159200 48282 160000 6 IRQ[2]
port 114 nsew signal input
rlabel metal2 s 79138 159200 79194 160000 6 IRQ[3]
port 115 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 IRQ[4]
port 116 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 IRQ[5]
port 117 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 IRQ[6]
port 118 nsew signal input
rlabel metal2 s 106922 159200 106978 160000 6 IRQ[7]
port 119 nsew signal input
rlabel metal2 s 110050 159200 110106 160000 6 IRQ[8]
port 120 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 IRQ[9]
port 121 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 NMI
port 122 nsew signal input
rlabel metal3 s 119200 122408 120000 122528 6 SYSTICKCLKDIV[0]
port 123 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 SYSTICKCLKDIV[10]
port 124 nsew signal input
rlabel metal3 s 119200 154504 120000 154624 6 SYSTICKCLKDIV[11]
port 125 nsew signal input
rlabel metal3 s 119200 117784 120000 117904 6 SYSTICKCLKDIV[12]
port 126 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 SYSTICKCLKDIV[13]
port 127 nsew signal input
rlabel metal2 s 23386 159200 23442 160000 6 SYSTICKCLKDIV[14]
port 128 nsew signal input
rlabel metal2 s 103794 159200 103850 160000 6 SYSTICKCLKDIV[15]
port 129 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 SYSTICKCLKDIV[16]
port 130 nsew signal input
rlabel metal2 s 57426 159200 57482 160000 6 SYSTICKCLKDIV[17]
port 131 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 SYSTICKCLKDIV[18]
port 132 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 SYSTICKCLKDIV[19]
port 133 nsew signal input
rlabel metal3 s 119200 94936 120000 95056 6 SYSTICKCLKDIV[1]
port 134 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 SYSTICKCLKDIV[20]
port 135 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 SYSTICKCLKDIV[21]
port 136 nsew signal input
rlabel metal2 s 41970 159200 42026 160000 6 SYSTICKCLKDIV[22]
port 137 nsew signal input
rlabel metal3 s 119200 76712 120000 76832 6 SYSTICKCLKDIV[23]
port 138 nsew signal input
rlabel metal3 s 119200 99560 120000 99680 6 SYSTICKCLKDIV[2]
port 139 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 SYSTICKCLKDIV[3]
port 140 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 SYSTICKCLKDIV[4]
port 141 nsew signal input
rlabel metal3 s 119200 145256 120000 145376 6 SYSTICKCLKDIV[5]
port 142 nsew signal input
rlabel metal2 s 32586 159200 32642 160000 6 SYSTICKCLKDIV[6]
port 143 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 SYSTICKCLKDIV[7]
port 144 nsew signal input
rlabel metal2 s 113178 159200 113234 160000 6 SYSTICKCLKDIV[8]
port 145 nsew signal input
rlabel metal2 s 60554 159200 60610 160000 6 SYSTICKCLKDIV[9]
port 146 nsew signal input
rlabel metal4 s 96368 2128 96688 157808 6 VPWR
port 147 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 VPWR
port 148 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 VPWR
port 149 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 150 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 VGND
port 151 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 VGND
port 152 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 VGND
port 153 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 VGND
port 154 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 120000 160000
string LEFview TRUE
<< end >>
