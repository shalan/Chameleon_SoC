magic
tech sky130A
magscale 1 2
timestamp 1608831475
<< obsli1 >>
rect 1104 2159 119019 77809
<< obsm1 >>
rect 474 892 119494 79144
<< metal2 >>
rect 754 79200 810 80000
rect 2226 79200 2282 80000
rect 3698 79200 3754 80000
rect 5170 79200 5226 80000
rect 6734 79200 6790 80000
rect 8206 79200 8262 80000
rect 9678 79200 9734 80000
rect 11242 79200 11298 80000
rect 12714 79200 12770 80000
rect 14186 79200 14242 80000
rect 15750 79200 15806 80000
rect 17222 79200 17278 80000
rect 18694 79200 18750 80000
rect 20166 79200 20222 80000
rect 21730 79200 21786 80000
rect 23202 79200 23258 80000
rect 24674 79200 24730 80000
rect 26238 79200 26294 80000
rect 27710 79200 27766 80000
rect 29182 79200 29238 80000
rect 30746 79200 30802 80000
rect 32218 79200 32274 80000
rect 33690 79200 33746 80000
rect 35162 79200 35218 80000
rect 36726 79200 36782 80000
rect 38198 79200 38254 80000
rect 39670 79200 39726 80000
rect 41234 79200 41290 80000
rect 42706 79200 42762 80000
rect 44178 79200 44234 80000
rect 45742 79200 45798 80000
rect 47214 79200 47270 80000
rect 48686 79200 48742 80000
rect 50158 79200 50214 80000
rect 51722 79200 51778 80000
rect 53194 79200 53250 80000
rect 54666 79200 54722 80000
rect 56230 79200 56286 80000
rect 57702 79200 57758 80000
rect 59174 79200 59230 80000
rect 60738 79200 60794 80000
rect 62210 79200 62266 80000
rect 63682 79200 63738 80000
rect 65154 79200 65210 80000
rect 66718 79200 66774 80000
rect 68190 79200 68246 80000
rect 69662 79200 69718 80000
rect 71226 79200 71282 80000
rect 72698 79200 72754 80000
rect 74170 79200 74226 80000
rect 75734 79200 75790 80000
rect 77206 79200 77262 80000
rect 78678 79200 78734 80000
rect 80150 79200 80206 80000
rect 81714 79200 81770 80000
rect 83186 79200 83242 80000
rect 84658 79200 84714 80000
rect 86222 79200 86278 80000
rect 87694 79200 87750 80000
rect 89166 79200 89222 80000
rect 90730 79200 90786 80000
rect 92202 79200 92258 80000
rect 93674 79200 93730 80000
rect 95146 79200 95202 80000
rect 96710 79200 96766 80000
rect 98182 79200 98238 80000
rect 99654 79200 99710 80000
rect 101218 79200 101274 80000
rect 102690 79200 102746 80000
rect 104162 79200 104218 80000
rect 105726 79200 105782 80000
rect 107198 79200 107254 80000
rect 108670 79200 108726 80000
rect 110142 79200 110198 80000
rect 111706 79200 111762 80000
rect 113178 79200 113234 80000
rect 114650 79200 114706 80000
rect 116214 79200 116270 80000
rect 117686 79200 117742 80000
rect 119158 79200 119214 80000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11702 0 11758 800
rect 12622 0 12678 800
rect 13542 0 13598 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17314 0 17370 800
rect 18234 0 18290 800
rect 19154 0 19210 800
rect 20074 0 20130 800
rect 21086 0 21142 800
rect 22006 0 22062 800
rect 22926 0 22982 800
rect 23846 0 23902 800
rect 24766 0 24822 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32310 0 32366 800
rect 33230 0 33286 800
rect 34150 0 34206 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38842 0 38898 800
rect 39762 0 39818 800
rect 40774 0 40830 800
rect 41694 0 41750 800
rect 42614 0 42670 800
rect 43534 0 43590 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46386 0 46442 800
rect 47306 0 47362 800
rect 48226 0 48282 800
rect 49146 0 49202 800
rect 50066 0 50122 800
rect 51078 0 51134 800
rect 51998 0 52054 800
rect 52918 0 52974 800
rect 53838 0 53894 800
rect 54758 0 54814 800
rect 55770 0 55826 800
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58530 0 58586 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61382 0 61438 800
rect 62302 0 62358 800
rect 63222 0 63278 800
rect 64142 0 64198 800
rect 65062 0 65118 800
rect 66074 0 66130 800
rect 66994 0 67050 800
rect 67914 0 67970 800
rect 68834 0 68890 800
rect 69754 0 69810 800
rect 70766 0 70822 800
rect 71686 0 71742 800
rect 72606 0 72662 800
rect 73526 0 73582 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 78218 0 78274 800
rect 79138 0 79194 800
rect 80058 0 80114 800
rect 81070 0 81126 800
rect 81990 0 82046 800
rect 82910 0 82966 800
rect 83830 0 83886 800
rect 84750 0 84806 800
rect 85762 0 85818 800
rect 86682 0 86738 800
rect 87602 0 87658 800
rect 88522 0 88578 800
rect 89442 0 89498 800
rect 90454 0 90510 800
rect 91374 0 91430 800
rect 92294 0 92350 800
rect 93214 0 93270 800
rect 94134 0 94190 800
rect 95054 0 95110 800
rect 96066 0 96122 800
rect 96986 0 97042 800
rect 97906 0 97962 800
rect 98826 0 98882 800
rect 99746 0 99802 800
rect 100758 0 100814 800
rect 101678 0 101734 800
rect 102598 0 102654 800
rect 103518 0 103574 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106370 0 106426 800
rect 107290 0 107346 800
rect 108210 0 108266 800
rect 109130 0 109186 800
rect 110050 0 110106 800
rect 111062 0 111118 800
rect 111982 0 112038 800
rect 112902 0 112958 800
rect 113822 0 113878 800
rect 114742 0 114798 800
rect 115754 0 115810 800
rect 116674 0 116730 800
rect 117594 0 117650 800
rect 118514 0 118570 800
rect 119434 0 119490 800
<< obsm2 >>
rect 480 79144 698 79200
rect 866 79144 2170 79200
rect 2338 79144 3642 79200
rect 3810 79144 5114 79200
rect 5282 79144 6678 79200
rect 6846 79144 8150 79200
rect 8318 79144 9622 79200
rect 9790 79144 11186 79200
rect 11354 79144 12658 79200
rect 12826 79144 14130 79200
rect 14298 79144 15694 79200
rect 15862 79144 17166 79200
rect 17334 79144 18638 79200
rect 18806 79144 20110 79200
rect 20278 79144 21674 79200
rect 21842 79144 23146 79200
rect 23314 79144 24618 79200
rect 24786 79144 26182 79200
rect 26350 79144 27654 79200
rect 27822 79144 29126 79200
rect 29294 79144 30690 79200
rect 30858 79144 32162 79200
rect 32330 79144 33634 79200
rect 33802 79144 35106 79200
rect 35274 79144 36670 79200
rect 36838 79144 38142 79200
rect 38310 79144 39614 79200
rect 39782 79144 41178 79200
rect 41346 79144 42650 79200
rect 42818 79144 44122 79200
rect 44290 79144 45686 79200
rect 45854 79144 47158 79200
rect 47326 79144 48630 79200
rect 48798 79144 50102 79200
rect 50270 79144 51666 79200
rect 51834 79144 53138 79200
rect 53306 79144 54610 79200
rect 54778 79144 56174 79200
rect 56342 79144 57646 79200
rect 57814 79144 59118 79200
rect 59286 79144 60682 79200
rect 60850 79144 62154 79200
rect 62322 79144 63626 79200
rect 63794 79144 65098 79200
rect 65266 79144 66662 79200
rect 66830 79144 68134 79200
rect 68302 79144 69606 79200
rect 69774 79144 71170 79200
rect 71338 79144 72642 79200
rect 72810 79144 74114 79200
rect 74282 79144 75678 79200
rect 75846 79144 77150 79200
rect 77318 79144 78622 79200
rect 78790 79144 80094 79200
rect 80262 79144 81658 79200
rect 81826 79144 83130 79200
rect 83298 79144 84602 79200
rect 84770 79144 86166 79200
rect 86334 79144 87638 79200
rect 87806 79144 89110 79200
rect 89278 79144 90674 79200
rect 90842 79144 92146 79200
rect 92314 79144 93618 79200
rect 93786 79144 95090 79200
rect 95258 79144 96654 79200
rect 96822 79144 98126 79200
rect 98294 79144 99598 79200
rect 99766 79144 101162 79200
rect 101330 79144 102634 79200
rect 102802 79144 104106 79200
rect 104274 79144 105670 79200
rect 105838 79144 107142 79200
rect 107310 79144 108614 79200
rect 108782 79144 110086 79200
rect 110254 79144 111650 79200
rect 111818 79144 113122 79200
rect 113290 79144 114594 79200
rect 114762 79144 116158 79200
rect 116326 79144 117630 79200
rect 117798 79144 119102 79200
rect 119270 79144 119488 79200
rect 480 856 119488 79144
rect 590 800 1342 856
rect 1510 800 2262 856
rect 2430 800 3182 856
rect 3350 800 4102 856
rect 4270 800 5022 856
rect 5190 800 6034 856
rect 6202 800 6954 856
rect 7122 800 7874 856
rect 8042 800 8794 856
rect 8962 800 9714 856
rect 9882 800 10726 856
rect 10894 800 11646 856
rect 11814 800 12566 856
rect 12734 800 13486 856
rect 13654 800 14406 856
rect 14574 800 15418 856
rect 15586 800 16338 856
rect 16506 800 17258 856
rect 17426 800 18178 856
rect 18346 800 19098 856
rect 19266 800 20018 856
rect 20186 800 21030 856
rect 21198 800 21950 856
rect 22118 800 22870 856
rect 23038 800 23790 856
rect 23958 800 24710 856
rect 24878 800 25722 856
rect 25890 800 26642 856
rect 26810 800 27562 856
rect 27730 800 28482 856
rect 28650 800 29402 856
rect 29570 800 30414 856
rect 30582 800 31334 856
rect 31502 800 32254 856
rect 32422 800 33174 856
rect 33342 800 34094 856
rect 34262 800 35014 856
rect 35182 800 36026 856
rect 36194 800 36946 856
rect 37114 800 37866 856
rect 38034 800 38786 856
rect 38954 800 39706 856
rect 39874 800 40718 856
rect 40886 800 41638 856
rect 41806 800 42558 856
rect 42726 800 43478 856
rect 43646 800 44398 856
rect 44566 800 45410 856
rect 45578 800 46330 856
rect 46498 800 47250 856
rect 47418 800 48170 856
rect 48338 800 49090 856
rect 49258 800 50010 856
rect 50178 800 51022 856
rect 51190 800 51942 856
rect 52110 800 52862 856
rect 53030 800 53782 856
rect 53950 800 54702 856
rect 54870 800 55714 856
rect 55882 800 56634 856
rect 56802 800 57554 856
rect 57722 800 58474 856
rect 58642 800 59394 856
rect 59562 800 60406 856
rect 60574 800 61326 856
rect 61494 800 62246 856
rect 62414 800 63166 856
rect 63334 800 64086 856
rect 64254 800 65006 856
rect 65174 800 66018 856
rect 66186 800 66938 856
rect 67106 800 67858 856
rect 68026 800 68778 856
rect 68946 800 69698 856
rect 69866 800 70710 856
rect 70878 800 71630 856
rect 71798 800 72550 856
rect 72718 800 73470 856
rect 73638 800 74390 856
rect 74558 800 75402 856
rect 75570 800 76322 856
rect 76490 800 77242 856
rect 77410 800 78162 856
rect 78330 800 79082 856
rect 79250 800 80002 856
rect 80170 800 81014 856
rect 81182 800 81934 856
rect 82102 800 82854 856
rect 83022 800 83774 856
rect 83942 800 84694 856
rect 84862 800 85706 856
rect 85874 800 86626 856
rect 86794 800 87546 856
rect 87714 800 88466 856
rect 88634 800 89386 856
rect 89554 800 90398 856
rect 90566 800 91318 856
rect 91486 800 92238 856
rect 92406 800 93158 856
rect 93326 800 94078 856
rect 94246 800 94998 856
rect 95166 800 96010 856
rect 96178 800 96930 856
rect 97098 800 97850 856
rect 98018 800 98770 856
rect 98938 800 99690 856
rect 99858 800 100702 856
rect 100870 800 101622 856
rect 101790 800 102542 856
rect 102710 800 103462 856
rect 103630 800 104382 856
rect 104550 800 105394 856
rect 105562 800 106314 856
rect 106482 800 107234 856
rect 107402 800 108154 856
rect 108322 800 109074 856
rect 109242 800 109994 856
rect 110162 800 111006 856
rect 111174 800 111926 856
rect 112094 800 112846 856
rect 113014 800 113766 856
rect 113934 800 114686 856
rect 114854 800 115698 856
rect 115866 800 116618 856
rect 116786 800 117538 856
rect 117706 800 118458 856
rect 118626 800 119378 856
<< metal3 >>
rect 0 69912 800 70032
rect 0 49920 800 50040
rect 0 29928 800 30048
rect 0 9936 800 10056
<< obsm3 >>
rect 800 70112 118207 77825
rect 880 69832 118207 70112
rect 800 50120 118207 69832
rect 880 49840 118207 50120
rect 800 30128 118207 49840
rect 880 29848 118207 30128
rect 800 10136 118207 29848
rect 880 9856 118207 10136
rect 800 2143 118207 9856
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
rect 81008 2128 81328 77840
rect 96368 2128 96688 77840
rect 111728 2128 112048 77840
<< obsm4 >>
rect 21955 3979 34848 75309
rect 35328 3979 50208 75309
rect 50688 3979 65568 75309
rect 66048 3979 80928 75309
rect 81408 3979 96288 75309
rect 96768 3979 109973 75309
<< labels >>
rlabel metal2 s 754 79200 810 80000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 15750 79200 15806 80000 6 A[10]
port 2 nsew signal input
rlabel metal2 s 17222 79200 17278 80000 6 A[11]
port 3 nsew signal input
rlabel metal2 s 18694 79200 18750 80000 6 A[12]
port 4 nsew signal input
rlabel metal2 s 20166 79200 20222 80000 6 A[13]
port 5 nsew signal input
rlabel metal2 s 21730 79200 21786 80000 6 A[14]
port 6 nsew signal input
rlabel metal2 s 23202 79200 23258 80000 6 A[15]
port 7 nsew signal input
rlabel metal2 s 24674 79200 24730 80000 6 A[16]
port 8 nsew signal input
rlabel metal2 s 26238 79200 26294 80000 6 A[17]
port 9 nsew signal input
rlabel metal2 s 27710 79200 27766 80000 6 A[18]
port 10 nsew signal input
rlabel metal2 s 29182 79200 29238 80000 6 A[19]
port 11 nsew signal input
rlabel metal2 s 2226 79200 2282 80000 6 A[1]
port 12 nsew signal input
rlabel metal2 s 30746 79200 30802 80000 6 A[20]
port 13 nsew signal input
rlabel metal2 s 32218 79200 32274 80000 6 A[21]
port 14 nsew signal input
rlabel metal2 s 33690 79200 33746 80000 6 A[22]
port 15 nsew signal input
rlabel metal2 s 35162 79200 35218 80000 6 A[23]
port 16 nsew signal input
rlabel metal2 s 3698 79200 3754 80000 6 A[2]
port 17 nsew signal input
rlabel metal2 s 5170 79200 5226 80000 6 A[3]
port 18 nsew signal input
rlabel metal2 s 6734 79200 6790 80000 6 A[4]
port 19 nsew signal input
rlabel metal2 s 8206 79200 8262 80000 6 A[5]
port 20 nsew signal input
rlabel metal2 s 9678 79200 9734 80000 6 A[6]
port 21 nsew signal input
rlabel metal2 s 11242 79200 11298 80000 6 A[7]
port 22 nsew signal input
rlabel metal2 s 12714 79200 12770 80000 6 A[8]
port 23 nsew signal input
rlabel metal2 s 14186 79200 14242 80000 6 A[9]
port 24 nsew signal input
rlabel metal2 s 36726 79200 36782 80000 6 A_h[0]
port 25 nsew signal input
rlabel metal2 s 51722 79200 51778 80000 6 A_h[10]
port 26 nsew signal input
rlabel metal2 s 53194 79200 53250 80000 6 A_h[11]
port 27 nsew signal input
rlabel metal2 s 54666 79200 54722 80000 6 A_h[12]
port 28 nsew signal input
rlabel metal2 s 56230 79200 56286 80000 6 A_h[13]
port 29 nsew signal input
rlabel metal2 s 57702 79200 57758 80000 6 A_h[14]
port 30 nsew signal input
rlabel metal2 s 59174 79200 59230 80000 6 A_h[15]
port 31 nsew signal input
rlabel metal2 s 60738 79200 60794 80000 6 A_h[16]
port 32 nsew signal input
rlabel metal2 s 62210 79200 62266 80000 6 A_h[17]
port 33 nsew signal input
rlabel metal2 s 63682 79200 63738 80000 6 A_h[18]
port 34 nsew signal input
rlabel metal2 s 65154 79200 65210 80000 6 A_h[19]
port 35 nsew signal input
rlabel metal2 s 38198 79200 38254 80000 6 A_h[1]
port 36 nsew signal input
rlabel metal2 s 66718 79200 66774 80000 6 A_h[20]
port 37 nsew signal input
rlabel metal2 s 68190 79200 68246 80000 6 A_h[21]
port 38 nsew signal input
rlabel metal2 s 69662 79200 69718 80000 6 A_h[22]
port 39 nsew signal input
rlabel metal2 s 71226 79200 71282 80000 6 A_h[23]
port 40 nsew signal input
rlabel metal2 s 39670 79200 39726 80000 6 A_h[2]
port 41 nsew signal input
rlabel metal2 s 41234 79200 41290 80000 6 A_h[3]
port 42 nsew signal input
rlabel metal2 s 42706 79200 42762 80000 6 A_h[4]
port 43 nsew signal input
rlabel metal2 s 44178 79200 44234 80000 6 A_h[5]
port 44 nsew signal input
rlabel metal2 s 45742 79200 45798 80000 6 A_h[6]
port 45 nsew signal input
rlabel metal2 s 47214 79200 47270 80000 6 A_h[7]
port 46 nsew signal input
rlabel metal2 s 48686 79200 48742 80000 6 A_h[8]
port 47 nsew signal input
rlabel metal2 s 50158 79200 50214 80000 6 A_h[9]
port 48 nsew signal input
rlabel metal2 s 72698 79200 72754 80000 6 Do[0]
port 49 nsew signal output
rlabel metal2 s 87694 79200 87750 80000 6 Do[10]
port 50 nsew signal output
rlabel metal2 s 89166 79200 89222 80000 6 Do[11]
port 51 nsew signal output
rlabel metal2 s 90730 79200 90786 80000 6 Do[12]
port 52 nsew signal output
rlabel metal2 s 92202 79200 92258 80000 6 Do[13]
port 53 nsew signal output
rlabel metal2 s 93674 79200 93730 80000 6 Do[14]
port 54 nsew signal output
rlabel metal2 s 95146 79200 95202 80000 6 Do[15]
port 55 nsew signal output
rlabel metal2 s 96710 79200 96766 80000 6 Do[16]
port 56 nsew signal output
rlabel metal2 s 98182 79200 98238 80000 6 Do[17]
port 57 nsew signal output
rlabel metal2 s 99654 79200 99710 80000 6 Do[18]
port 58 nsew signal output
rlabel metal2 s 101218 79200 101274 80000 6 Do[19]
port 59 nsew signal output
rlabel metal2 s 74170 79200 74226 80000 6 Do[1]
port 60 nsew signal output
rlabel metal2 s 102690 79200 102746 80000 6 Do[20]
port 61 nsew signal output
rlabel metal2 s 104162 79200 104218 80000 6 Do[21]
port 62 nsew signal output
rlabel metal2 s 105726 79200 105782 80000 6 Do[22]
port 63 nsew signal output
rlabel metal2 s 107198 79200 107254 80000 6 Do[23]
port 64 nsew signal output
rlabel metal2 s 108670 79200 108726 80000 6 Do[24]
port 65 nsew signal output
rlabel metal2 s 110142 79200 110198 80000 6 Do[25]
port 66 nsew signal output
rlabel metal2 s 111706 79200 111762 80000 6 Do[26]
port 67 nsew signal output
rlabel metal2 s 113178 79200 113234 80000 6 Do[27]
port 68 nsew signal output
rlabel metal2 s 114650 79200 114706 80000 6 Do[28]
port 69 nsew signal output
rlabel metal2 s 116214 79200 116270 80000 6 Do[29]
port 70 nsew signal output
rlabel metal2 s 75734 79200 75790 80000 6 Do[2]
port 71 nsew signal output
rlabel metal2 s 117686 79200 117742 80000 6 Do[30]
port 72 nsew signal output
rlabel metal2 s 119158 79200 119214 80000 6 Do[31]
port 73 nsew signal output
rlabel metal2 s 77206 79200 77262 80000 6 Do[3]
port 74 nsew signal output
rlabel metal2 s 78678 79200 78734 80000 6 Do[4]
port 75 nsew signal output
rlabel metal2 s 80150 79200 80206 80000 6 Do[5]
port 76 nsew signal output
rlabel metal2 s 81714 79200 81770 80000 6 Do[6]
port 77 nsew signal output
rlabel metal2 s 83186 79200 83242 80000 6 Do[7]
port 78 nsew signal output
rlabel metal2 s 84658 79200 84714 80000 6 Do[8]
port 79 nsew signal output
rlabel metal2 s 86222 79200 86278 80000 6 Do[9]
port 80 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 clk
port 81 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 hit
port 82 nsew signal output
rlabel metal2 s 478 0 534 800 6 line[0]
port 83 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 line[100]
port 84 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 line[101]
port 85 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 line[102]
port 86 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 line[103]
port 87 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 line[104]
port 88 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 line[105]
port 89 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 line[106]
port 90 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 line[107]
port 91 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 line[108]
port 92 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 line[109]
port 93 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 line[10]
port 94 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 line[110]
port 95 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 line[111]
port 96 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 line[112]
port 97 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 line[113]
port 98 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 line[114]
port 99 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 line[115]
port 100 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 line[116]
port 101 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 line[117]
port 102 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 line[118]
port 103 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 line[119]
port 104 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 line[11]
port 105 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 line[120]
port 106 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 line[121]
port 107 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 line[122]
port 108 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 line[123]
port 109 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 line[124]
port 110 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 line[125]
port 111 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 line[126]
port 112 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 line[127]
port 113 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 line[12]
port 114 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 line[13]
port 115 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 line[14]
port 116 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 line[15]
port 117 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 line[16]
port 118 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 line[17]
port 119 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 line[18]
port 120 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 line[19]
port 121 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 line[1]
port 122 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 line[20]
port 123 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 line[21]
port 124 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 line[22]
port 125 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 line[23]
port 126 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 line[24]
port 127 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 line[25]
port 128 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 line[26]
port 129 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 line[27]
port 130 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 line[28]
port 131 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 line[29]
port 132 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 line[2]
port 133 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 line[30]
port 134 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 line[31]
port 135 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 line[32]
port 136 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 line[33]
port 137 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 line[34]
port 138 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 line[35]
port 139 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 line[36]
port 140 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 line[37]
port 141 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 line[38]
port 142 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 line[39]
port 143 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 line[3]
port 144 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 line[40]
port 145 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 line[41]
port 146 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 line[42]
port 147 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 line[43]
port 148 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 line[44]
port 149 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 line[45]
port 150 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 line[46]
port 151 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 line[47]
port 152 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 line[48]
port 153 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 line[49]
port 154 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 line[4]
port 155 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 line[50]
port 156 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 line[51]
port 157 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 line[52]
port 158 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 line[53]
port 159 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 line[54]
port 160 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 line[55]
port 161 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 line[56]
port 162 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 line[57]
port 163 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 line[58]
port 164 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 line[59]
port 165 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 line[5]
port 166 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 line[60]
port 167 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 line[61]
port 168 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 line[62]
port 169 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 line[63]
port 170 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 line[64]
port 171 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 line[65]
port 172 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 line[66]
port 173 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 line[67]
port 174 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 line[68]
port 175 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 line[69]
port 176 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 line[6]
port 177 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 line[70]
port 178 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 line[71]
port 179 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 line[72]
port 180 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 line[73]
port 181 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 line[74]
port 182 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 line[75]
port 183 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 line[76]
port 184 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 line[77]
port 185 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 line[78]
port 186 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 line[79]
port 187 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 line[7]
port 188 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 line[80]
port 189 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 line[81]
port 190 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 line[82]
port 191 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 line[83]
port 192 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 line[84]
port 193 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 line[85]
port 194 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 line[86]
port 195 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 line[87]
port 196 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 line[88]
port 197 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 line[89]
port 198 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 line[8]
port 199 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 line[90]
port 200 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 line[91]
port 201 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 line[92]
port 202 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 line[93]
port 203 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 line[94]
port 204 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 line[95]
port 205 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 line[96]
port 206 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 line[97]
port 207 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 line[98]
port 208 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 line[99]
port 209 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 line[9]
port 210 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rst_n
port 211 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 wr
port 212 nsew signal input
rlabel metal4 s 96368 2128 96688 77840 6 VPWR
port 213 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 VPWR
port 214 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 VPWR
port 215 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 77840 6 VPWR
port 216 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 77840 6 VGND
port 217 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 77840 6 VGND
port 218 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 VGND
port 219 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 VGND
port 220 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 119494 80000
string LEFview TRUE
<< end >>
