* NGSPICE file created from DMC_32x16HC.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

.subckt DMC_32x16HC A[0] A[10] A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19]
+ A[1] A[20] A[21] A[22] A[23] A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A_h[0] A_h[10]
+ A_h[11] A_h[12] A_h[13] A_h[14] A_h[15] A_h[16] A_h[17] A_h[18] A_h[19] A_h[1] A_h[20]
+ A_h[21] A_h[22] A_h[23] A_h[2] A_h[3] A_h[4] A_h[5] A_h[6] A_h[7] A_h[8] A_h[9]
+ Do[0] Do[10] Do[11] Do[12] Do[13] Do[14] Do[15] Do[16] Do[17] Do[18] Do[19] Do[1]
+ Do[20] Do[21] Do[22] Do[23] Do[24] Do[25] Do[26] Do[27] Do[28] Do[29] Do[2] Do[30]
+ Do[31] Do[3] Do[4] Do[5] Do[6] Do[7] Do[8] Do[9] clk hit line[0] line[100] line[101]
+ line[102] line[103] line[104] line[105] line[106] line[107] line[108] line[109]
+ line[10] line[110] line[111] line[112] line[113] line[114] line[115] line[116] line[117]
+ line[118] line[119] line[11] line[120] line[121] line[122] line[123] line[124] line[125]
+ line[126] line[127] line[12] line[13] line[14] line[15] line[16] line[17] line[18]
+ line[19] line[1] line[20] line[21] line[22] line[23] line[24] line[25] line[26]
+ line[27] line[28] line[29] line[2] line[30] line[31] line[32] line[33] line[34]
+ line[35] line[36] line[37] line[38] line[39] line[3] line[40] line[41] line[42]
+ line[43] line[44] line[45] line[46] line[47] line[48] line[49] line[4] line[50]
+ line[51] line[52] line[53] line[54] line[55] line[56] line[57] line[58] line[59]
+ line[5] line[60] line[61] line[62] line[63] line[64] line[65] line[66] line[67]
+ line[68] line[69] line[6] line[70] line[71] line[72] line[73] line[74] line[75]
+ line[76] line[77] line[78] line[79] line[7] line[80] line[81] line[82] line[83]
+ line[84] line[85] line[86] line[87] line[88] line[89] line[8] line[90] line[91]
+ line[92] line[93] line[94] line[95] line[96] line[97] line[98] line[99] line[9]
+ rst_n wr VPWR VGND
XOVHB\[16\].VALID\[10\].TOBUF OVHB\[16\].VALID\[10\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09515__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05903_ _05903_/A _05922_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_06883_ _06883_/A _06902_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_09671_ _09670_/Q _09702_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05834_ _05836_/CLK line[18] VGND VGND VPWR VPWR _05835_/A sky130_fd_sc_hd__dfxtp_1
X_08622_ _08646_/CLK line[27] VGND VGND VPWR VPWR _08622_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ _08552_/Q _08582_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05765_ _05764_/Q _05782_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11780__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06874__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07504_ _07518_/CLK line[28] VGND VGND VPWR VPWR _07504_/Q sky130_fd_sc_hd__dfxtp_1
X_08484_ _08480_/CLK line[92] VGND VGND VPWR VPWR _08485_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05696_ _05708_/CLK line[83] VGND VGND VPWR VPWR _05697_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09250__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10396__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07435_ _07434_/Q _07462_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07366_ _07380_/CLK line[93] VGND VGND VPWR VPWR _07367_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09105_ _09105_/CLK _09106_/X VGND VGND VPWR VPWR _09085_/CLK sky130_fd_sc_hd__dlclkp_1
X_06317_ _06317_/A _06342_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_07297_ _07296_/Q _07322_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_09036_ _13923_/X wr VGND VGND VPWR VPWR _09036_/X sky130_fd_sc_hd__and2_1
X_06248_ _06244_/CLK line[94] VGND VGND VPWR VPWR _06248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[27\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06179_ _06179_/A _06202_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11020__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06114__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11955__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04929__A1_N A_h[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09938_ _09937_/Q _09947_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05953__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09425__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06411__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09869_ _09849_/CLK line[71] VGND VGND VPWR VPWR _09869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11900_ _11900_/A _11907_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_12880_ _12879_/Q _12887_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_11831_ _11823_/CLK line[72] VGND VGND VPWR VPWR _11831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11762_ _11762_/A _11767_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13497_/CLK line[67] VGND VGND VPWR VPWR _13501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10707_/CLK line[73] VGND VGND VPWR VPWR _10713_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11691_/CLK line[9] VGND VGND VPWR VPWR _11693_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13431_/Q _13447_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10644_ _10644_/A _10647_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10575_ _10575_/CLK _10576_/X VGND VGND VPWR VPWR _10571_/CLK sky130_fd_sc_hd__dlclkp_1
X_13363_ _13347_/CLK line[4] VGND VGND VPWR VPWR _13363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12314_ _12313_/Q _12327_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08504__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13294_ _13293_/Q _13307_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_12245_ _12227_/CLK line[5] VGND VGND VPWR VPWR _12246_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12176_ _12176_/A _12187_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_11127_ _11111_/CLK line[6] VGND VGND VPWR VPWR _11127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[0\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05863__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11058_ _11057_/Q _11067_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10009_ _10011_/CLK line[7] VGND VGND VPWR VPWR _10009_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12696__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].CGAND _13923_/X wr VGND VGND VPWR VPWR OVHB\[22\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_45_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05550_ _05568_/CLK line[31] VGND VGND VPWR VPWR _05550_/Q sky130_fd_sc_hd__dfxtp_1
X_05481_ _05480_/Q _05502_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11105__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07220_ _07232_/CLK line[26] VGND VGND VPWR VPWR _07221_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05103__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07151_ _07150_/Q _07182_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10944__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13320__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06102_ _06108_/CLK line[27] VGND VGND VPWR VPWR _06103_/A sky130_fd_sc_hd__dfxtp_1
X_07082_ _07098_/CLK line[91] VGND VGND VPWR VPWR _07082_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08414__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06033_ _06032_/Q _06062_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[1\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[4\].TOBUF OVHB\[18\].VALID\[4\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07984_ _07983_/Q _07987_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09723_ _09721_/CLK line[4] VGND VGND VPWR VPWR _09723_/Q sky130_fd_sc_hd__dfxtp_1
X_06935_ _06935_/CLK _06936_/X VGND VGND VPWR VPWR _06923_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_41_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13990__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09654_ _09653_/Q _09667_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06866_ _06832_/A wr VGND VGND VPWR VPWR _06866_/X sky130_fd_sc_hd__and2_1
X_08605_ _08609_/CLK line[5] VGND VGND VPWR VPWR _08606_/A sky130_fd_sc_hd__dfxtp_1
X_05817_ _13910_/X VGND VGND VPWR VPWR _05817_/Y sky130_fd_sc_hd__inv_2
X_09585_ _09577_/CLK line[69] VGND VGND VPWR VPWR _09585_/Q sky130_fd_sc_hd__dfxtp_1
X_06797_ _06832_/A VGND VGND VPWR VPWR _06797_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08536_ _08535_/Q _08547_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_05748_ _05756_/CLK line[112] VGND VGND VPWR VPWR _05748_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _08473_/CLK line[70] VGND VGND VPWR VPWR _08468_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05679_ _05679_/A _05712_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ _07417_/Q _07427_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_08398_ _08397_/Q _08407_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05013__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ _07327_/CLK line[71] VGND VGND VPWR VPWR _07349_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[9\].FF OVHB\[9\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[9\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10360_ _10360_/A _10367_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_09019_ _09005_/CLK line[66] VGND VGND VPWR VPWR _09019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10291_ _10277_/CLK line[8] VGND VGND VPWR VPWR _10292_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12030_ _12029_/Q _12047_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11685__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06779__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09155__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13981_ A_h[5] VGND VGND VPWR VPWR _13990_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_DATA\[25\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[9\]_A0 _11414_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08994__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ _12931_/Q _12957_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[24\].VALID\[3\].TOBUF OVHB\[24\].VALID\[3\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12863_ _12881_/CLK line[46] VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11814_ _11813_/Q _11837_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12794_ _12793_/Q _12817_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07403__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11745_ _11757_/CLK line[47] VGND VGND VPWR VPWR _11746_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06019__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11676_ _11676_/A _11697_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05501__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13415_ _13439_/CLK line[42] VGND VGND VPWR VPWR _13415_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10627_ _10627_/CLK line[33] VGND VGND VPWR VPWR _10628_/A sky130_fd_sc_hd__dfxtp_1
X_13346_ _13346_/A _13377_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_10558_ _10557_/Q _10577_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13277_ _13285_/CLK line[107] VGND VGND VPWR VPWR _13277_/Q sky130_fd_sc_hd__dfxtp_1
X_10489_ _10473_/CLK line[98] VGND VGND VPWR VPWR _10489_/Q sky130_fd_sc_hd__dfxtp_1
X_12228_ _12228_/A _12257_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[24\]_A3 _12777_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11595__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12159_ _12177_/CLK line[108] VGND VGND VPWR VPWR _12159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05593__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04981_ _04980_/Q _05012_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06720_ _06719_/Q _06727_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06651_ _06633_/CLK line[8] VGND VGND VPWR VPWR _06651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05602_ _05602_/A _05607_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_09370_ _09370_/A _09387_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
X_06582_ _06581_/Q _06587_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[9\].TOBUF OVHB\[16\].VALID\[9\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_08321_ _08329_/CLK line[3] VGND VGND VPWR VPWR _08321_/Q sky130_fd_sc_hd__dfxtp_1
X_05533_ _05519_/CLK line[9] VGND VGND VPWR VPWR _05533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ _08251_/Q _08267_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_05464_ _05463_/Q _05467_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[2\].TOBUF OVHB\[30\].VALID\[2\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_07203_ _07183_/CLK line[4] VGND VGND VPWR VPWR _07203_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10674__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08183_ _08175_/CLK line[68] VGND VGND VPWR VPWR _08184_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05395_ _05395_/CLK _05396_/X VGND VGND VPWR VPWR _05391_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13050__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05768__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07134_ _07133_/Q _07147_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08144__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08722__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[1\].FF OVHB\[18\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[18\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13985__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07065_ _07043_/CLK line[69] VGND VGND VPWR VPWR _07066_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07983__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08441__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06016_ _06016_/A _06027_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[12\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07967_ _07981_/CLK line[97] VGND VGND VPWR VPWR _07967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].CGAND_A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09706_ _09705_/Q _09737_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06918_ _06918_/A _06937_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07898_ _07898_/A _07917_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05008__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09703__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09637_ _09659_/CLK line[107] VGND VGND VPWR VPWR _09638_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10849__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06849_ _06839_/CLK line[98] VGND VGND VPWR VPWR _06850_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13225__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08319__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09568_ _09567_/Q _09597_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08519_ _08541_/CLK line[108] VGND VGND VPWR VPWR _08519_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _09507_/CLK line[44] VGND VGND VPWR VPWR _09499_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[27\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _11530_/A _11557_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10584__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11461_ _11479_/CLK line[45] VGND VGND VPWR VPWR _11462_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05678__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13200_ _13200_/CLK _13201_/X VGND VGND VPWR VPWR _13194_/CLK sky130_fd_sc_hd__dlclkp_1
X_10412_ _10411_/Q _10437_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
X_11392_ _11391_/Q _11417_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[8\].TOBUF OVHB\[22\].VALID\[8\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _13272_/A wr VGND VGND VPWR VPWR _13131_/X sky130_fd_sc_hd__and2_1
X_10343_ _10341_/CLK line[46] VGND VGND VPWR VPWR _10343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07893__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10274_ _10273_/Q _10297_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_13062_ _12992_/A VGND VGND VPWR VPWR _13062_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12013_ _12019_/CLK line[32] VGND VGND VPWR VPWR _12013_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[12\].TOBUF OVHB\[6\].VALID\[12\].FF/Q OVHB\[6\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_79_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[16\].VALID\[3\].FF OVHB\[16\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[16\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05991__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13964_ _13960_/X _13964_/B _13958_/X _13966_/D VGND VGND VPWR VPWR _13964_/X sky130_fd_sc_hd__and4b_4
XANTENNA__10402__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10759__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12915_ _12914_/Q _12922_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10121__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13895_ _13894_/Q _13902_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13135__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12846_ _12820_/CLK line[24] VGND VGND VPWR VPWR _12846_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07133__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[23\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12974__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12777_ _12776_/Q _12782_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11728_ _11706_/CLK line[25] VGND VGND VPWR VPWR _11728_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11659_ _11658_/Q _11662_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05180_ _05179_/Q _05187_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[16\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13329_ _13328_/Q _13342_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06062__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12214__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08870_ _08869_/Q _08897_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07308__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07821_ _07837_/CLK line[45] VGND VGND VPWR VPWR _07822_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07752_ _07751_/Q _07777_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_04964_ _04963_/Q _04977_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09523__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06703_ _06711_/CLK line[46] VGND VGND VPWR VPWR _06704_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[0\].TOBUF OVHB\[6\].VALID\[0\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[26\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07683_ _07679_/CLK line[110] VGND VGND VPWR VPWR _07684_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ _09352_/A VGND VGND VPWR VPWR _09422_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06634_ _06633_/Q _06657_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[5\].FF OVHB\[14\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[14\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07043__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09353_ _09365_/CLK line[96] VGND VGND VPWR VPWR _09353_/Q sky130_fd_sc_hd__dfxtp_1
X_06565_ _06565_/CLK line[111] VGND VGND VPWR VPWR _06566_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[9\].FF OVHB\[31\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[31\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08304_ _08303_/Q _08337_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_05516_ _05515_/Q _05537_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06882__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09284_ _09283_/Q _09317_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_06496_ _06495_/Q _06517_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06237__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05447_ _05445_/CLK line[97] VGND VGND VPWR VPWR _05448_/A sky130_fd_sc_hd__dfxtp_1
X_08235_ _08257_/CLK line[106] VGND VGND VPWR VPWR _08235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05498__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05378_ _05378_/A _05397_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_08166_ _08165_/Q _08197_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ _07117_/CLK line[107] VGND VGND VPWR VPWR _07117_/Q sky130_fd_sc_hd__dfxtp_1
X_08097_ _08113_/CLK line[43] VGND VGND VPWR VPWR _08098_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07048_ _07047_/Q _07077_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12124__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07218__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06122__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08999_ _08999_/A _09002_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11963__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[29\].VALID\[14\].TOBUF OVHB\[29\].VALID\[14\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__04935__B2 _04935_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09433__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10961_ _11032_/A wr VGND VGND VPWR VPWR _10961_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.MUX\[6\]_A3 _13578_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12700_ _12708_/CLK line[85] VGND VGND VPWR VPWR _12700_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08049__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13680_ _13682_/CLK line[21] VGND VGND VPWR VPWR _13681_/A sky130_fd_sc_hd__dfxtp_1
X_10892_ _11032_/A VGND VGND VPWR VPWR _10892_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07531__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12631_ _12630_/Q _12642_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[14\]_A2 _13494_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12560_/CLK line[22] VGND VGND VPWR VPWR _12562_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _11512_/Q _11522_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12492_/Q _12502_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10892__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[24\].INV _13972_/Y VGND VGND VPWR VPWR OVHB\[24\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__11203__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[12\].VALID\[7\].FF OVHB\[12\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[12\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11444_ _11440_/CLK line[23] VGND VGND VPWR VPWR _11445_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11375_ _11375_/A _11382_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09608__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13114_ _13120_/CLK line[18] VGND VGND VPWR VPWR _13114_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[13\].TOBUF OVHB\[22\].VALID\[13\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10326_ _10314_/CLK line[24] VGND VGND VPWR VPWR _10326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13045_ _13045_/A _13062_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_10257_ _10257_/A _10262_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].V OVHB\[24\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[24\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06032__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07706__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10188_ _10188_/CLK line[89] VGND VGND VPWR VPWR _10189_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11873__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05871__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10489__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13947_ A_h[4] VGND VGND VPWR VPWR _13950_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13878_ _13882_/CLK line[126] VGND VGND VPWR VPWR _13879_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10786__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12829_ _12828_/Q _12852_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07798__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06350_ _06349_/Q _06377_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05301_ _05299_/CLK line[45] VGND VGND VPWR VPWR _05301_/Q sky130_fd_sc_hd__dfxtp_1
X_06281_ _06285_/CLK line[109] VGND VGND VPWR VPWR _06281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[29\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _10960_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11113__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05232_ _05231_/Q _05257_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_08020_ _08020_/CLK _08021_/X VGND VGND VPWR VPWR _08000_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06207__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05111__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10952__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05163_ _05157_/CLK line[110] VGND VGND VPWR VPWR _05163_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[5\].TOBUF OVHB\[4\].VALID\[5\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_6_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[10\].VOBUF OVHB\[10\].V/Q OVHB\[10\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__08422__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09971_ _09970_/Q _09982_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_05094_ _05093_/Q _05117_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[29\].VALID\[8\].TOBUF OVHB\[29\].VALID\[8\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_08922_ _08922_/CLK line[22] VGND VGND VPWR VPWR _08923_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[9\].FF OVHB\[10\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[10\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].V OVHB\[15\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[15\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07038__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12879__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08853_ _08852_/Q _08862_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[30\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07804_ _07788_/CLK line[23] VGND VGND VPWR VPWR _07804_/Q sky130_fd_sc_hd__dfxtp_1
X_08784_ _08762_/CLK line[87] VGND VGND VPWR VPWR _08784_/Q sky130_fd_sc_hd__dfxtp_1
X_05996_ _05995_/Q _06027_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07735_ _07735_/A _07742_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_04947_ _04947_/CLK line[11] VGND VGND VPWR VPWR _04947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07666_ _07644_/CLK line[88] VGND VGND VPWR VPWR _07666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[23\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09405_ _09405_/A _09422_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_06617_ _06616_/Q _06622_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_07597_ _07596_/Q _07602_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13503__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09336_ _09320_/CLK line[83] VGND VGND VPWR VPWR _09336_/Q sky130_fd_sc_hd__dfxtp_1
X_06548_ _06528_/CLK line[89] VGND VGND VPWR VPWR _06549_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09267_ _09267_/A _09282_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_06479_ _06478_/Q _06482_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_08218_ _08208_/CLK line[84] VGND VGND VPWR VPWR _08219_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05021__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09198_ _09200_/CLK line[20] VGND VGND VPWR VPWR _09198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10862__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08149_ _08148_/Q _08162_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[28\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _10575_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11160_ _11148_/CLK line[21] VGND VGND VPWR VPWR _11160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10111_ _10110_/Q _10122_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_11091_ _11090_/Q _11102_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12432__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[18\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _07705_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10042_ _10042_/CLK line[22] VGND VGND VPWR VPWR _10042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12789__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11693__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12151__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06787__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09163__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[0\].TOBUF OVHB\[11\].VALID\[0\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05046__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13801_ _13800_/Q _13832_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11993_ _11992_/Q _12012_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10102__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13732_ _13746_/CLK line[59] VGND VGND VPWR VPWR _13733_/A sky130_fd_sc_hd__dfxtp_1
X_10944_ _10930_/CLK line[50] VGND VGND VPWR VPWR _10944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ _13662_/Q _13692_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_10875_ _10874_/Q _10892_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13413__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ _12638_/CLK line[60] VGND VGND VPWR VPWR _12614_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ _13598_/CLK line[124] VGND VGND VPWR VPWR _13594_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07411__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12029__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12545_ _12545_/A _12572_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12607__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12476_ _12490_/CLK line[125] VGND VGND VPWR VPWR _12476_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08092__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11868__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12326__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[0\].FF OVHB\[5\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[5\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11427_ _11426_/Q _11452_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[18\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[16\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09338__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11358_ _11370_/CLK line[126] VGND VGND VPWR VPWR _11358_/Q sky130_fd_sc_hd__dfxtp_1
X_10309_ _10308_/Q _10332_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_11289_ _11288_/Q _11312_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_13028_ _13050_/CLK line[112] VGND VGND VPWR VPWR _13028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06697__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05850_ _05850_/CLK _05851_/X VGND VGND VPWR VPWR _05836_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09073__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _07320_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_94_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05781_ _13909_/X wr VGND VGND VPWR VPWR _05781_/X sky130_fd_sc_hd__and2_1
X_07520_ _07518_/CLK line[21] VGND VGND VPWR VPWR _07520_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09801__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08267__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07451_ _07451_/A _07462_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13901__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06402_ _06408_/CLK line[22] VGND VGND VPWR VPWR _06402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__04945__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07382_ _07380_/CLK line[86] VGND VGND VPWR VPWR _07382_/Q sky130_fd_sc_hd__dfxtp_1
X_09121_ _09120_/Q _09142_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_06333_ _06332_/Q _06342_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09052_ _09068_/CLK line[81] VGND VGND VPWR VPWR _09053_/A sky130_fd_sc_hd__dfxtp_1
X_06264_ _06244_/CLK line[87] VGND VGND VPWR VPWR _06265_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11778__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08003_ _08003_/A _08022_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_05215_ _05215_/A _05222_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_06195_ _06194_/Q _06202_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09248__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05776__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05146_ _05122_/CLK line[88] VGND VGND VPWR VPWR _05146_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08152__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].CGAND _13918_/X wr VGND VGND VPWR VPWR OVHB\[17\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05077_ _05076_/Q _05082_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_09954_ _09978_/CLK line[124] VGND VGND VPWR VPWR _09954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08905_ _08904_/Q _08932_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[2\].FF OVHB\[3\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[3\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09885_ _09884_/Q _09912_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08836_ _08850_/CLK line[125] VGND VGND VPWR VPWR _08837_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12402__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09561__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06400__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08767_ _08766_/Q _08792_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05979_ _05978_/Q _05992_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11018__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07718_ _07724_/CLK line[126] VGND VGND VPWR VPWR _07719_/A sky130_fd_sc_hd__dfxtp_1
X_08698_ _08710_/CLK line[62] VGND VGND VPWR VPWR _08699_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09711__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07649_ _07649_/A _07672_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[16\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _06935_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13233__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10660_ _10656_/CLK line[63] VGND VGND VPWR VPWR _10660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08327__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[9\].INV _13951_/X VGND VGND VPWR VPWR OVHB\[9\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09319_ _09318_/Q _09352_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_10591_ _10591_/A _10612_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_12330_ _12352_/CLK line[58] VGND VGND VPWR VPWR _12330_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10592__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12261_ _12260_/Q _12292_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05686__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11212_ _11216_/CLK line[59] VGND VGND VPWR VPWR _11212_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08062__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09736__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _12204_/CLK line[123] VGND VGND VPWR VPWR _12193_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11143_ _11142_/Q _11172_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_11074_ _11090_/CLK line[124] VGND VGND VPWR VPWR _11074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13408__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[12\].TOBUF OVHB\[19\].VALID\[12\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10025_ _10024_/Q _10052_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06310__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11976_ _12151_/A wr VGND VGND VPWR VPWR _11976_/X sky130_fd_sc_hd__and2_1
XFILLER_91_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[1\].VALID\[4\].FF OVHB\[1\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[1\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13715_ _13701_/CLK line[37] VGND VGND VPWR VPWR _13715_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10767__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10927_ _11032_/A VGND VGND VPWR VPWR _10927_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13143__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08237__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XMUX.MUX\[8\] _09452_/Z _10922_/Z _10992_/Z _13582_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[8] sky130_fd_sc_hd__mux4_1
X_13646_ _13645_/Q _13657_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_10858_ _10872_/CLK line[16] VGND VGND VPWR VPWR _10858_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07141__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12982__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13577_ _13559_/CLK line[102] VGND VGND VPWR VPWR _13577_/Q sky130_fd_sc_hd__dfxtp_1
X_10789_ _10788_/Q _10822_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11241__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12528_ _12528_/A _12537_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12459_ _12449_/CLK line[103] VGND VGND VPWR VPWR _12459_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[11\].TOBUF OVHB\[12\].VALID\[11\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09068__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05000_ _05000_/CLK line[21] VGND VGND VPWR VPWR _05000_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[27\]_A1 _10373_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10007__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08700__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06951_ _06950_/Q _06972_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[14\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13318__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05902_ _05902_/CLK line[49] VGND VGND VPWR VPWR _05903_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _09694_/CLK line[122] VGND VGND VPWR VPWR _09670_/Q sky130_fd_sc_hd__dfxtp_1
X_06882_ _06892_/CLK line[113] VGND VGND VPWR VPWR _06883_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07316__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08621_ _08620_/Q _08652_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_05833_ _05832_/Q _05852_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11416__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08552_ _08560_/CLK line[123] VGND VGND VPWR VPWR _08552_/Q sky130_fd_sc_hd__dfxtp_1
X_05764_ _05756_/CLK line[114] VGND VGND VPWR VPWR _05764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[18\].VALID\[0\].TOBUF OVHB\[18\].VALID\[0\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_07503_ _07503_/A _07532_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_08483_ _08482_/Q _08512_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05695_ _05694_/Q _05712_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_07434_ _07446_/CLK line[124] VGND VGND VPWR VPWR _07434_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07051__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13988__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12892__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07365_ _07364_/Q _07392_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_09104_ _09104_/A _09107_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_06316_ _06320_/CLK line[125] VGND VGND VPWR VPWR _06317_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06890__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[7\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07296_ _07292_/CLK line[61] VGND VGND VPWR VPWR _07296_/Q sky130_fd_sc_hd__dfxtp_1
X_09035_ _09035_/CLK _09036_/X VGND VGND VPWR VPWR _09005_/CLK sky130_fd_sc_hd__dlclkp_1
X_06247_ _06246_/Q _06272_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06178_ _06186_/CLK line[62] VGND VGND VPWR VPWR _06179_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05129_ _05128_/Q _05152_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07076__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09937_ _09925_/CLK line[102] VGND VGND VPWR VPWR _09937_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12132__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09868_ _09867_/Q _09877_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07226__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08819_ _08823_/CLK line[103] VGND VGND VPWR VPWR _08819_/Q sky130_fd_sc_hd__dfxtp_1
X_09799_ _09793_/CLK line[39] VGND VGND VPWR VPWR _09799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11971__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11830_ _11829_/Q _11837_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09441__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11761_ _11757_/CLK line[40] VGND VGND VPWR VPWR _11762_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13499_/Q _13517_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10711_/Q _10717_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11692_/A _11697_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13898__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13431_ _13439_/CLK line[35] VGND VGND VPWR VPWR _13431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10643_ _10627_/CLK line[41] VGND VGND VPWR VPWR _10644_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13362_ _13361_/Q _13377_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10574_ _10573_/Q _10577_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12313_ _12311_/CLK line[36] VGND VGND VPWR VPWR _12313_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12307__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13293_ _13285_/CLK line[100] VGND VGND VPWR VPWR _13293_/Q sky130_fd_sc_hd__dfxtp_1
X_12244_ _12243_/Q _12257_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_12175_ _12177_/CLK line[101] VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09616__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11126_ _11126_/A _11137_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11057_ _11063_/CLK line[102] VGND VGND VPWR VPWR _11057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06040__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10008_ _10007_/Q _10017_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[24\].VALID\[14\].FF OVHB\[24\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[24\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11881__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06975__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10497__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11959_ _11945_/CLK line[2] VGND VGND VPWR VPWR _11959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[3\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05480_ _05476_/CLK line[127] VGND VGND VPWR VPWR _05480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[26\].VALID\[1\].FF OVHB\[26\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[26\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13629_ _13631_/CLK line[12] VGND VGND VPWR VPWR _13629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ _07170_/CLK line[122] VGND VGND VPWR VPWR _07150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06101_ _06100_/Q _06132_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_07081_ _07081_/A _07112_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11121__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06032_ _06050_/CLK line[123] VGND VGND VPWR VPWR _06032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06215__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[5\].TOBUF OVHB\[16\].VALID\[5\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08430__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07983_ _07981_/CLK line[105] VGND VGND VPWR VPWR _07983_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13048__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09722_ _09722_/A _09737_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_06934_ _06933_/Q _06937_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[8\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _13620_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_83_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09653_ _09659_/CLK line[100] VGND VGND VPWR VPWR _09653_/Q sky130_fd_sc_hd__dfxtp_1
X_06865_ _06865_/CLK _06866_/X VGND VGND VPWR VPWR _06839_/CLK sky130_fd_sc_hd__dlclkp_1
X_08604_ _08604_/A _08617_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05816_ _13910_/X wr VGND VGND VPWR VPWR _05816_/X sky130_fd_sc_hd__and2_1
X_09584_ _09583_/Q _09597_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_06796_ _06832_/A wr VGND VGND VPWR VPWR _06796_/X sky130_fd_sc_hd__and2_1
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08535_ _08541_/CLK line[101] VGND VGND VPWR VPWR _08535_/Q sky130_fd_sc_hd__dfxtp_1
X_05747_ _13909_/X VGND VGND VPWR VPWR _05747_/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[12\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _08465_/Q _08477_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05678_ _05708_/CLK line[80] VGND VGND VPWR VPWR _05679_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _07393_/CLK line[102] VGND VGND VPWR VPWR _07417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _08383_/CLK line[38] VGND VGND VPWR VPWR _08397_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13511__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07348_ _07348_/A _07357_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08605__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07279_ _07267_/CLK line[39] VGND VGND VPWR VPWR _07279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[24\].VALID\[3\].FF OVHB\[24\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[24\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09018_ _09018_/A _09037_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10290_ _10290_/A _10297_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10870__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05964__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08340__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13980_ A_h[4] VGND VGND VPWR VPWR _13990_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_MUX.MUX\[9\]_A1 _12884_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[31\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12931_ _12937_/CLK line[77] VGND VGND VPWR VPWR _12931_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12797__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[22\].VALID\[4\].TOBUF OVHB\[22\].VALID\[4\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_12862_ _12861_/Q _12887_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[7\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _13235_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09171__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11813_ _11823_/CLK line[78] VGND VGND VPWR VPWR _11813_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[17\]_A0 _10873_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ _12803_/CLK line[14] VGND VGND VPWR VPWR _12793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13271__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10110__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11744_ _11743_/Q _11767_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05204__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11675_ _11691_/CLK line[15] VGND VGND VPWR VPWR _11676_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13421__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13413_/Q _13447_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08515__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10626_ _10625_/Q _10647_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05501__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12037__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13345_ _13347_/CLK line[10] VGND VGND VPWR VPWR _13346_/A sky130_fd_sc_hd__dfxtp_1
X_10557_ _10571_/CLK line[1] VGND VGND VPWR VPWR _10557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13276_ _13275_/Q _13307_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_10488_ _10487_/Q _10507_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12227_ _12227_/CLK line[11] VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09346__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12158_ _12158_/A _12187_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13446__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11109_ _11111_/CLK line[12] VGND VGND VPWR VPWR _11109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12089_ _12109_/CLK line[76] VGND VGND VPWR VPWR _12089_/Q sky130_fd_sc_hd__dfxtp_1
X_04980_ _05000_/CLK line[26] VGND VGND VPWR VPWR _04980_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[5\].FF OVHB\[22\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[22\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[10\].FF OVHB\[30\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[30\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06650_ _06650_/A _06657_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09081__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05601_ _05575_/CLK line[40] VGND VGND VPWR VPWR _05602_/A sky130_fd_sc_hd__dfxtp_1
X_06581_ _06565_/CLK line[104] VGND VGND VPWR VPWR _06581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _08319_/Q _08337_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10020__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05532_ _05531_/Q _05537_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08251_ _08257_/CLK line[99] VGND VGND VPWR VPWR _08251_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[6\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _12850_/CLK sky130_fd_sc_hd__clkbuf_4
X_05463_ _05445_/CLK line[105] VGND VGND VPWR VPWR _05463_/Q sky130_fd_sc_hd__dfxtp_1
X_07202_ _07201_/Q _07217_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04953__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08182_ _08181_/Q _08197_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_05394_ _05394_/A _05397_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07133_ _07117_/CLK line[100] VGND VGND VPWR VPWR _07133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07064_ _07063_/Q _07077_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11786__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06015_ _06023_/CLK line[101] VGND VGND VPWR VPWR _06016_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[12\].FF OVHB\[20\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[20\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09256__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[9\].VALID\[14\].TOBUF OVHB\[9\].VALID\[14\].FF/Q OVHB\[9\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_102_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07966_ _07965_/Q _07987_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[16\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09705_ _09721_/CLK line[10] VGND VGND VPWR VPWR _09705_/Q sky130_fd_sc_hd__dfxtp_1
X_06917_ _06923_/CLK line[1] VGND VGND VPWR VPWR _06918_/A sky130_fd_sc_hd__dfxtp_1
X_07897_ _07905_/CLK line[65] VGND VGND VPWR VPWR _07898_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09636_ _09635_/Q _09667_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12410__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06848_ _06847_/Q _06867_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _10190_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07504__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09567_ _09577_/CLK line[75] VGND VGND VPWR VPWR _09567_/Q sky130_fd_sc_hd__dfxtp_1
X_06779_ _06775_/CLK line[66] VGND VGND VPWR VPWR _06779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11026__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[20\].VALID\[7\].FF OVHB\[20\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[20\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08518_ _08517_/Q _08547_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _09497_/Q _09527_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _08473_/CLK line[76] VGND VGND VPWR VPWR _08449_/Q sky130_fd_sc_hd__dfxtp_1
XMUX.MUX\[26\] _11421_/Z _13451_/Z _06521_/Z _13591_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[26] sky130_fd_sc_hd__mux4_1
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[10\].VALID\[14\].FF OVHB\[10\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[10\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ _11460_/A _11487_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VALID\[10\].TOBUF OVHB\[29\].VALID\[10\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[10\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10411_ _10405_/CLK line[77] VGND VGND VPWR VPWR _10411_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[13\].TOBUF OVHB\[2\].VALID\[13\].FF/Q OVHB\[2\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_11391_ _11395_/CLK line[13] VGND VGND VPWR VPWR _11391_/Q sky130_fd_sc_hd__dfxtp_1
X_13130_ _13130_/CLK _13131_/X VGND VGND VPWR VPWR _13120_/CLK sky130_fd_sc_hd__dlclkp_1
X_10342_ _10341_/Q _10367_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[9\].TOBUF OVHB\[20\].VALID\[9\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_13061_ _12992_/A wr VGND VGND VPWR VPWR _13061_/X sky130_fd_sc_hd__and2_1
X_10273_ _10277_/CLK line[14] VGND VGND VPWR VPWR _10273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05694__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ _12151_/A VGND VGND VPWR VPWR _12012_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08070__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05991__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13963_ _13960_/X _13958_/X _13964_/B _13966_/D VGND VGND VPWR VPWR _13963_/X sky130_fd_sc_hd__and4bb_4
XFILLER_101_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[3\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12914_ _12902_/CLK line[55] VGND VGND VPWR VPWR _12914_/Q sky130_fd_sc_hd__dfxtp_1
X_13894_ _13882_/CLK line[119] VGND VGND VPWR VPWR _13894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[8\].FF OVHB\[19\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[19\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12845_ _12845_/A _12852_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_12776_ _12774_/CLK line[120] VGND VGND VPWR VPWR _12776_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[25\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _09805_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10775__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11727_ _11727_/A _11732_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13151__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05869__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08245__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11658_ _11636_/CLK line[121] VGND VGND VPWR VPWR _11658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _10608_/Q _10612_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11589_ _11589_/A _11592_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_13328_ _13308_/CLK line[116] VGND VGND VPWR VPWR _13328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[11\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13259_ _13258_/Q _13272_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07820_ _07819_/Q _07847_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05109__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07751_ _07773_/CLK line[13] VGND VGND VPWR VPWR _07751_/Q sky130_fd_sc_hd__dfxtp_1
X_04963_ _04947_/CLK line[4] VGND VGND VPWR VPWR _04963_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13326__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06702_ _06701_/Q _06727_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13904__A A[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07682_ _07681_/Q _07707_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_09421_ _09352_/A wr VGND VGND VPWR VPWR _09421_/X sky130_fd_sc_hd__and2_1
X_06633_ _06633_/CLK line[14] VGND VGND VPWR VPWR _06633_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[1\].TOBUF OVHB\[4\].VALID\[1\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_09352_ _09352_/A VGND VGND VPWR VPWR _09352_/Y sky130_fd_sc_hd__inv_2
XOVHB\[29\].VALID\[4\].TOBUF OVHB\[29\].VALID\[4\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_06564_ _06564_/A _06587_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08303_ _08329_/CLK line[0] VGND VGND VPWR VPWR _08303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10685__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05515_ _05519_/CLK line[15] VGND VGND VPWR VPWR _05515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09283_ _09307_/CLK line[64] VGND VGND VPWR VPWR _09283_/Q sky130_fd_sc_hd__dfxtp_1
X_06495_ _06489_/CLK line[79] VGND VGND VPWR VPWR _06495_/Q sky130_fd_sc_hd__dfxtp_1
X_08234_ _08233_/Q _08267_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_05446_ _05445_/Q _05467_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_08165_ _08175_/CLK line[74] VGND VGND VPWR VPWR _08165_/Q sky130_fd_sc_hd__dfxtp_1
X_05377_ _05391_/CLK line[65] VGND VGND VPWR VPWR _05378_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07994__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07116_ _07116_/A _07147_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08096_ _08095_/Q _08127_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[14\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _06550_/CLK sky130_fd_sc_hd__clkbuf_4
X_07047_ _07043_/CLK line[75] VGND VGND VPWR VPWR _07047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08998_ _08972_/CLK line[57] VGND VGND VPWR VPWR _08999_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05019__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07949_ _07948_/Q _07952_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[31\].CGAND_A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12140__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10960_ _10960_/CLK _10961_/X VGND VGND VPWR VPWR _10930_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07234__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07812__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09619_ _09618_/Q _09632_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10891_ _11032_/A wr VGND VGND VPWR VPWR _10891_/X sky130_fd_sc_hd__and2_1
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _12638_/CLK line[53] VGND VGND VPWR VPWR _12630_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[22\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07531__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[14\]_A3 _05164_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12560_/Q _12572_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[24\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _11500_/CLK line[54] VGND VGND VPWR VPWR _11512_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12490_/CLK line[118] VGND VGND VPWR VPWR _12492_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11443_ _11442_/Q _11452_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[30\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11374_ _11370_/CLK line[119] VGND VGND VPWR VPWR _11375_/A sky130_fd_sc_hd__dfxtp_1
X_13113_ _13112_/Q _13132_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12315__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10325_ _10325_/A _10332_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07409__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[14\].FF OVHB\[29\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[29\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13044_ _13050_/CLK line[114] VGND VGND VPWR VPWR _13045_/A sky130_fd_sc_hd__dfxtp_1
X_10256_ _10248_/CLK line[120] VGND VGND VPWR VPWR _10257_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07706__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[13\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _06165_/CLK sky130_fd_sc_hd__clkbuf_4
X_10187_ _10186_/Q _10192_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09624__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12050__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13946_ _13944_/B _13946_/B _13944_/C _13944_/D VGND VGND VPWR VPWR _13272_/A sky130_fd_sc_hd__and4_4
XFILLER_62_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[12\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ _13876_/Q _13902_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06983__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12828_ _12820_/CLK line[30] VGND VGND VPWR VPWR _12828_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A _12782_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].CG clk OVHB\[4\].CGAND/X VGND VGND VPWR VPWR OVHB\[4\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05599__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05300_ _05300_/A _05327_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_06280_ _06279_/Q _06307_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_05231_ _05253_/CLK line[13] VGND VGND VPWR VPWR _05231_/Q sky130_fd_sc_hd__dfxtp_1
X_05162_ _05162_/A _05187_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12225__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09970_ _09978_/CLK line[117] VGND VGND VPWR VPWR _09970_/Q sky130_fd_sc_hd__dfxtp_1
X_05093_ _05093_/CLK line[78] VGND VGND VPWR VPWR _05093_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[6\].TOBUF OVHB\[2\].VALID\[6\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__06223__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08921_ _08920_/Q _08932_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[9\].TOBUF OVHB\[27\].VALID\[9\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08852_ _08850_/CLK line[118] VGND VGND VPWR VPWR _08852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09534__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07803_ _07802_/Q _07812_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_08783_ _08783_/A _08792_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_05995_ _06023_/CLK line[106] VGND VGND VPWR VPWR _05995_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13056__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07734_ _07724_/CLK line[119] VGND VGND VPWR VPWR _07735_/A sky130_fd_sc_hd__dfxtp_1
X_04946_ _04946_/A _04977_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_07665_ _07665_/A _07672_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09404_ _09414_/CLK line[114] VGND VGND VPWR VPWR _09405_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].CGAND _06272_/A wr VGND VGND VPWR VPWR OVHB\[13\].CG/GATE sky130_fd_sc_hd__and2_4
X_06616_ _06596_/CLK line[120] VGND VGND VPWR VPWR _06616_/Q sky130_fd_sc_hd__dfxtp_1
X_07596_ _07572_/CLK line[56] VGND VGND VPWR VPWR _07596_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05152__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09335_ _09334_/Q _09352_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_06547_ _06546_/Q _06552_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11304__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09266_ _09256_/CLK line[51] VGND VGND VPWR VPWR _09267_/A sky130_fd_sc_hd__dfxtp_1
X_06478_ _06464_/CLK line[57] VGND VGND VPWR VPWR _06478_/Q sky130_fd_sc_hd__dfxtp_1
X_08217_ _08216_/Q _08232_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05429_ _05428_/Q _05432_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_09197_ _09197_/A _09212_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09709__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08148_ _08134_/CLK line[52] VGND VGND VPWR VPWR _08148_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08613__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08079_ _08079_/A _08092_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10110_ _10100_/CLK line[53] VGND VGND VPWR VPWR _10110_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06133__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11090_ _11090_/CLK line[117] VGND VGND VPWR VPWR _11090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10041_ _10040_/Q _10052_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05972__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05327__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13800_ _13822_/CLK line[90] VGND VGND VPWR VPWR _13800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05046__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11992_ _12002_/CLK line[17] VGND VGND VPWR VPWR _11992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ _13730_/Q _13762_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_10943_ _10942_/Q _10962_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07899__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13662_ _13682_/CLK line[27] VGND VGND VPWR VPWR _13662_/Q sky130_fd_sc_hd__dfxtp_1
X_10874_ _10872_/CLK line[18] VGND VGND VPWR VPWR _10874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[1\].VALID\[14\].FF OVHB\[1\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[1\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ _12613_/A _12642_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13593_ _13592_/Q _13622_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11214__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06308__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12544_ _12560_/CLK line[28] VGND VGND VPWR VPWR _12545_/A sky130_fd_sc_hd__dfxtp_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05212__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12475_ _12474_/Q _12502_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[4\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08523__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11426_ _11440_/CLK line[29] VGND VGND VPWR VPWR _11426_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[22\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11357_ _11356_/Q _11382_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07139__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10308_ _10314_/CLK line[30] VGND VGND VPWR VPWR _10308_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06621__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11288_ _11302_/CLK line[94] VGND VGND VPWR VPWR _11288_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[5\].FF OVHB\[8\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[8\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13027_ _12992_/A VGND VGND VPWR VPWR _13027_/Y sky130_fd_sc_hd__inv_2
X_10239_ _10238_/Q _10262_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05780_ _05780_/CLK _05781_/X VGND VGND VPWR VPWR _05756_/CLK sky130_fd_sc_hd__dlclkp_1
X_13929_ _13934_/C _13934_/B _13933_/B _13934_/D VGND VGND VPWR VPWR _09912_/A sky130_fd_sc_hd__and4bb_4
XANTENNA__13604__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[27\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07450_ _07446_/CLK line[117] VGND VGND VPWR VPWR _07451_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06401_ _06400_/Q _06412_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13901__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07381_ _07381_/A _07392_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_09120_ _09116_/CLK line[127] VGND VGND VPWR VPWR _09120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06332_ _06320_/CLK line[118] VGND VGND VPWR VPWR _06332_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05122__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[12\].FF OVHB\[25\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[25\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10963__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09051_ _09050_/Q _09072_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_06263_ _06262_/Q _06272_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08002_ _08000_/CLK line[113] VGND VGND VPWR VPWR _08003_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04961__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05214_ _05214_/CLK line[119] VGND VGND VPWR VPWR _05215_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[4\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06194_ _06186_/CLK line[55] VGND VGND VPWR VPWR _06194_/Q sky130_fd_sc_hd__dfxtp_1
X_05145_ _05145_/A _05152_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07049__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05076_ _05058_/CLK line[56] VGND VGND VPWR VPWR _05076_/Q sky130_fd_sc_hd__dfxtp_1
X_09953_ _09952_/Q _09982_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11794__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06888__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08904_ _08922_/CLK line[28] VGND VGND VPWR VPWR _08904_/Q sky130_fd_sc_hd__dfxtp_1
X_09884_ _09908_/CLK line[92] VGND VGND VPWR VPWR _09884_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09264__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09842__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08835_ _08835_/A _08862_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VOBUF OVHB\[7\].V/Q OVHB\[7\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].INV _13968_/X VGND VGND VPWR VPWR OVHB\[23\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__10203__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09561__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08766_ _08762_/CLK line[93] VGND VGND VPWR VPWR _08766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05978_ _05984_/CLK line[84] VGND VGND VPWR VPWR _05978_/Q sky130_fd_sc_hd__dfxtp_1
X_07717_ _07717_/A _07742_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_04929_ A_h[12] _04927_/Y A_h[15] _04924_/Y VGND VGND VPWR VPWR _04929_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[15\].VALID\[14\].FF OVHB\[15\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[15\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[7\].FF OVHB\[6\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[6\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08697_ _08696_/Q _08722_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07648_ _07644_/CLK line[94] VGND VGND VPWR VPWR _07649_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07512__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07579_ _07578_/Q _07602_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09318_ _09320_/CLK line[80] VGND VGND VPWR VPWR _09318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06128__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10590_ _10594_/CLK line[31] VGND VGND VPWR VPWR _10591_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11969__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09249_ _09248_/Q _09282_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09439__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12260_ _12268_/CLK line[26] VGND VGND VPWR VPWR _12260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[15\].VALID\[13\].TOBUF OVHB\[15\].VALID\[13\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_11211_ _11210_/Q _11242_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09736__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12191_ _12190_/Q _12222_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11142_ _11148_/CLK line[27] VGND VGND VPWR VPWR _11142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06798__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11073_ _11073_/A _11102_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[6\].TOBUF OVHB\[9\].VALID\[6\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10024_ _10042_/CLK line[28] VGND VGND VPWR VPWR _10024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09902__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11975_ _11975_/CLK _11976_/X VGND VGND VPWR VPWR _11945_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_45_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13714_ _13713_/Q _13727_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10926_ _11032_/A wr VGND VGND VPWR VPWR _10926_/X sky130_fd_sc_hd__and2_1
X_13645_ _13631_/CLK line[5] VGND VGND VPWR VPWR _13645_/Q sky130_fd_sc_hd__dfxtp_1
X_10857_ _11032_/A VGND VGND VPWR VPWR _10857_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11522__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06038__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _13575_/Q _13587_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_10788_ _10804_/CLK line[112] VGND VGND VPWR VPWR _10788_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11879__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[4\].VALID\[9\].FF OVHB\[4\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[4\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11241__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10783__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12527_ _12523_/CLK line[6] VGND VGND VPWR VPWR _12528_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05877__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08253__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12458_ _12457_/Q _12467_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[27\]_A2 _11003_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11409_ _11395_/CLK line[7] VGND VGND VPWR VPWR _11409_/Q sky130_fd_sc_hd__dfxtp_1
X_12389_ _12387_/CLK line[71] VGND VGND VPWR VPWR _12389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[4\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _12465_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06950_ _06960_/CLK line[31] VGND VGND VPWR VPWR _06950_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05901_ _05900_/Q _05922_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06501__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[20\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06881_ _06880_/Q _06902_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11119__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08620_ _08646_/CLK line[26] VGND VGND VPWR VPWR _08620_/Q sky130_fd_sc_hd__dfxtp_1
X_05832_ _05836_/CLK line[17] VGND VGND VPWR VPWR _05832_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09812__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07182__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08551_ _08550_/Q _08582_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10958__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05763_ _05763_/A _05782_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11416__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13334__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07502_ _07518_/CLK line[27] VGND VGND VPWR VPWR _07503_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08428__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08482_ _08480_/CLK line[91] VGND VGND VPWR VPWR _08482_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[1\].TOBUF OVHB\[16\].VALID\[1\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_05694_ _05708_/CLK line[82] VGND VGND VPWR VPWR _05694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07433_ _07432_/Q _07462_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ _07380_/CLK line[92] VGND VGND VPWR VPWR _07364_/Q sky130_fd_sc_hd__dfxtp_1
X_09103_ _09085_/CLK line[105] VGND VGND VPWR VPWR _09104_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10693__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06315_ _06314_/Q _06342_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_07295_ _07294_/Q _07322_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05787__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09034_ _09033_/Q _09037_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08163__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06246_ _06244_/CLK line[93] VGND VGND VPWR VPWR _06246_/Q sky130_fd_sc_hd__dfxtp_1
X_06177_ _06177_/A _06202_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05128_ _05122_/CLK line[94] VGND VGND VPWR VPWR _05128_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07357__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13509__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09936_ _09935_/Q _09947_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_05059_ _05058_/Q _05082_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07076__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09867_ _09849_/CLK line[70] VGND VGND VPWR VPWR _09867_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[3\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _12080_/CLK sky130_fd_sc_hd__clkbuf_4
X_08818_ _08817_/Q _08827_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09798_ _09798_/A _09807_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05027__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10868__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08749_ _08749_/CLK line[71] VGND VGND VPWR VPWR _08749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13244__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[10\].FF OVHB\[21\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[21\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11760_ _11759_/Q _11767_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08338__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07242__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10711_ _10707_/CLK line[72] VGND VGND VPWR VPWR _10711_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11691_/CLK line[8] VGND VGND VPWR VPWR _11692_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _10642_/A _10647_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_13430_ _13429_/Q _13447_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13347_/CLK line[3] VGND VGND VPWR VPWR _13361_/Q sky130_fd_sc_hd__dfxtp_1
X_10573_ _10571_/CLK line[9] VGND VGND VPWR VPWR _10573_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09169__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12312_ _12311_/Q _12327_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[1\].FF OVHB\[13\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[13\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13292_ _13291_/Q _13307_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08651__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[0\].TOBUF OVHB\[22\].VALID\[0\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10108__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12243_ _12227_/CLK line[4] VGND VGND VPWR VPWR _12243_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[5\].FF OVHB\[30\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[30\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08801__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ _12173_/Q _12187_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[23\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _09420_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13419__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11125_ _11111_/CLK line[5] VGND VGND VPWR VPWR _11126_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12323__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[12\].FF OVHB\[11\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[11\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[19\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07417__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11056_ _11056_/A _11067_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10007_ _10011_/CLK line[6] VGND VGND VPWR VPWR _10007_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[2\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _11135_/CLK sky130_fd_sc_hd__clkbuf_4
X_11958_ _11957_/Q _11977_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07152__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08826__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12993__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10909_ _10903_/CLK line[34] VGND VGND VPWR VPWR _10909_/Q sky130_fd_sc_hd__dfxtp_1
X_11889_ _11901_/CLK line[98] VGND VGND VPWR VPWR _11890_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06991__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13628_ _13627_/Q _13657_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13559_ _13559_/CLK line[108] VGND VGND VPWR VPWR _13560_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09079__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06100_ _06108_/CLK line[26] VGND VGND VPWR VPWR _06100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07080_ _07098_/CLK line[90] VGND VGND VPWR VPWR _07081_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[6\].FF OVHB\[29\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[29\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05400__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06031_ _06031_/A _06062_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10018__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[6\].TOBUF OVHB\[14\].VALID\[6\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__12233__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07982_ _07982_/A _07987_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[3\].FF OVHB\[11\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[11\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07327__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[8\].INV _13950_/Y VGND VGND VPWR VPWR OVHB\[8\].INV/Y sky130_fd_sc_hd__inv_2
X_09721_ _09721_/CLK line[3] VGND VGND VPWR VPWR _09722_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06231__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06933_ _06923_/CLK line[9] VGND VGND VPWR VPWR _06933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[22\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _09035_/CLK sky130_fd_sc_hd__clkbuf_4
X_09652_ _09652_/A _09667_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_06864_ _06863_/Q _06867_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10331__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09542__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05815_ _05815_/CLK _05816_/X VGND VGND VPWR VPWR _05799_/CLK sky130_fd_sc_hd__dlclkp_1
X_08603_ _08609_/CLK line[4] VGND VGND VPWR VPWR _08604_/A sky130_fd_sc_hd__dfxtp_1
X_09583_ _09577_/CLK line[68] VGND VGND VPWR VPWR _09583_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06795_ _06795_/CLK _06796_/X VGND VGND VPWR VPWR _06775_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_103_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08534_ _08533_/Q _08547_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_05746_ _13909_/X wr VGND VGND VPWR VPWR _05746_/X sky130_fd_sc_hd__and2_1
XANTENNA__08158__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ _08473_/CLK line[69] VGND VGND VPWR VPWR _08465_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05677_ _13909_/X VGND VGND VPWR VPWR _05677_/Y sky130_fd_sc_hd__inv_2
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[9\].VALID\[10\].TOBUF OVHB\[9\].VALID\[10\].FF/Q OVHB\[9\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ _07415_/Q _07427_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ _08395_/Q _08407_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07347_ _07327_/CLK line[70] VGND VGND VPWR VPWR _07348_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12408__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06406__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07278_ _07277_/Q _07287_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09017_ _09005_/CLK line[65] VGND VGND VPWR VPWR _09018_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06229_ _06223_/CLK line[71] VGND VGND VPWR VPWR _06230_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10506__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09717__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[8\].FF OVHB\[27\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[27\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06141__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09919_ _09925_/CLK line[108] VGND VGND VPWR VPWR _09919_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11982__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[9\]_A2 _13514_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ _12929_/Q _12957_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[14\].FF OVHB\[6\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[6\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05980__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10598__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12881_/CLK line[45] VGND VGND VPWR VPWR _12861_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13552__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11812_ _11811_/Q _11837_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08068__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[5\].TOBUF OVHB\[20\].VALID\[5\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[17\]_A1 _07023_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[21\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _08650_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12792_ _12791_/Q _12817_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13271__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11743_ _11757_/CLK line[46] VGND VGND VPWR VPWR _11743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _05780_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06166__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11674_ _11673_/Q _11697_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13413_ _13439_/CLK line[32] VGND VGND VPWR VPWR _13413_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _10627_/CLK line[47] VGND VGND VPWR VPWR _10625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11222__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10556_ _10555_/Q _10577_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06316__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13344_ _13343_/Q _13377_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13275_ _13285_/CLK line[106] VGND VGND VPWR VPWR _13275_/Q sky130_fd_sc_hd__dfxtp_1
X_10487_ _10473_/CLK line[97] VGND VGND VPWR VPWR _10487_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08531__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12226_ _12225_/Q _12257_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13149__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13727__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12157_ _12177_/CLK line[107] VGND VGND VPWR VPWR _12158_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11108_ _11108_/A _11137_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12988__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13446__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12088_ _12087_/Q _12117_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11039_ _11063_/CLK line[108] VGND VGND VPWR VPWR _11040_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05890__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[17\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05600_ _05599_/Q _05607_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_06580_ _06579_/Q _06587_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05531_ _05519_/CLK line[8] VGND VGND VPWR VPWR _05531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13612__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08250_ _08249_/Q _08267_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08706__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05462_ _05462_/A _05467_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_07201_ _07183_/CLK line[3] VGND VGND VPWR VPWR _07201_/Q sky130_fd_sc_hd__dfxtp_1
X_08181_ _08175_/CLK line[67] VGND VGND VPWR VPWR _08181_/Q sky130_fd_sc_hd__dfxtp_1
X_05393_ _05391_/CLK line[73] VGND VGND VPWR VPWR _05394_/A sky130_fd_sc_hd__dfxtp_1
X_07132_ _07132_/A _07147_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09387__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _05395_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05130__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10971__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07063_ _07043_/CLK line[68] VGND VGND VPWR VPWR _07063_/Q sky130_fd_sc_hd__dfxtp_1
X_06014_ _06013_/Q _06027_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[29\].VALID\[0\].TOBUF OVHB\[29\].VALID\[0\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_134_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07057__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12898__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07965_ _07981_/CLK line[111] VGND VGND VPWR VPWR _07965_/Q sky130_fd_sc_hd__dfxtp_1
X_09704_ _09703_/Q _09737_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06916_ _06916_/A _06937_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06896__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09272__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07896_ _07895_/Q _07917_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ _09659_/CLK line[106] VGND VGND VPWR VPWR _09635_/Q sky130_fd_sc_hd__dfxtp_1
X_06847_ _06839_/CLK line[97] VGND VGND VPWR VPWR _06847_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10996__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10211__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06778_ _06778_/A _06797_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_09566_ _09565_/Q _09597_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05305__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[11\].TOBUF OVHB\[25\].VALID\[11\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05729_ _05739_/CLK line[98] VGND VGND VPWR VPWR _05729_/Q sky130_fd_sc_hd__dfxtp_1
X_08517_ _08541_/CLK line[107] VGND VGND VPWR VPWR _08517_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _09507_/CLK line[43] VGND VGND VPWR VPWR _09497_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13522__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08448_ _08447_/Q _08477_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12138__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08379_ _08383_/CLK line[44] VGND VGND VPWR VPWR _08380_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[19\] _10877_/Z _10387_/Z _07097_/Z _07167_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[19] sky130_fd_sc_hd__mux4_1
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10410_ _10409_/Q _10437_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11390_ _11390_/A _11417_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_10341_ _10341_/CLK line[45] VGND VGND VPWR VPWR _10341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09447__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13060_ _13060_/CLK _13061_/X VGND VGND VPWR VPWR _13050_/CLK sky130_fd_sc_hd__dlclkp_1
X_10272_ _10271_/Q _10297_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12011_ _12151_/A wr VGND VGND VPWR VPWR _12011_/X sky130_fd_sc_hd__and2_1
XFILLER_132_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__04938__B1 A_h[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11067__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12601__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13962_ _13960_/X _13964_/B _13958_/X _13966_/D VGND VGND VPWR VPWR _13962_/X sky130_fd_sc_hd__and4bb_4
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09182__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _12912_/Q _12922_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13893_ _13893_/A _13902_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_12844_ _12820_/CLK line[23] VGND VGND VPWR VPWR _12845_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12775_ _12774_/Q _12782_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_11726_ _11706_/CLK line[24] VGND VGND VPWR VPWR _11727_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07430__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[4\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12048__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11657_/A _11662_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06046__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10608_ _10594_/CLK line[25] VGND VGND VPWR VPWR _10608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11588_ _11588_/CLK line[89] VGND VGND VPWR VPWR _11589_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11887__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13327_ _13326_/Q _13342_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_10539_ _10538_/Q _10542_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09357__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08261__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[12\].FF OVHB\[2\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[2\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13258_ _13254_/CLK line[84] VGND VGND VPWR VPWR _13258_/Q sky130_fd_sc_hd__dfxtp_1
X_12209_ _12208_/Q _12222_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12361__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _13188_/Q _13202_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04929__B1 A_h[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12511__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07750_ _07749_/Q _07777_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_04962_ _04961_/Q _04977_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07605__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06701_ _06711_/CLK line[45] VGND VGND VPWR VPWR _06701_/Q sky130_fd_sc_hd__dfxtp_1
X_07681_ _07679_/CLK line[109] VGND VGND VPWR VPWR _07681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11127__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06632_ _06632_/A _06657_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09420_ _09420_/CLK _09421_/X VGND VGND VPWR VPWR _09414_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09820__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[2\].TOBUF OVHB\[2\].VALID\[2\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_06563_ _06565_/CLK line[110] VGND VGND VPWR VPWR _06564_/A sky130_fd_sc_hd__dfxtp_1
X_09351_ _09352_/A wr VGND VGND VPWR VPWR _09351_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[18\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[5\].TOBUF OVHB\[27\].VALID\[5\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_05514_ _05513_/Q _05537_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_08302_ _13940_/X VGND VGND VPWR VPWR _08302_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08436__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09282_ _09352_/A VGND VGND VPWR VPWR _09282_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06494_ _06493_/Q _06517_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08233_ _08257_/CLK line[96] VGND VGND VPWR VPWR _08233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05445_ _05445_/CLK line[111] VGND VGND VPWR VPWR _05445_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12536__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08164_ _08163_/Q _08197_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_05376_ _05375_/Q _05397_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[0\].FF OVHB\[0\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[0\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07115_ _07117_/CLK line[106] VGND VGND VPWR VPWR _07116_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[11\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08095_ _08113_/CLK line[42] VGND VGND VPWR VPWR _08095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05795__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08171__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07046_ _07046_/A _07077_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[26\].VALID\[10\].FF OVHB\[26\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[26\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08997_ _08996_/Q _09002_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07948_ _07946_/CLK line[89] VGND VGND VPWR VPWR _07948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07879_ _07879_/A _07882_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11037__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09618_ _09626_/CLK line[84] VGND VGND VPWR VPWR _09618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05035__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08196__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10890_ _10890_/CLK _10891_/X VGND VGND VPWR VPWR _10872_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.MUX\[22\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10876__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ _09549_/A _09562_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13252__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08346__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12560_ _12560_/CLK line[21] VGND VGND VPWR VPWR _12560_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[30\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _11510_/Q _11522_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12491_/A _12502_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ _11440_/CLK line[22] VGND VGND VPWR VPWR _11442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[16\].VALID\[12\].FF OVHB\[16\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[16\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11373_ _11372_/Q _11382_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11500__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13112_ _13120_/CLK line[17] VGND VGND VPWR VPWR _13112_/Q sky130_fd_sc_hd__dfxtp_1
X_10324_ _10314_/CLK line[23] VGND VGND VPWR VPWR _10325_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10116__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10255_ _10255_/A _10262_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_13043_ _13042_/Q _13062_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10186_ _10188_/CLK line[88] VGND VGND VPWR VPWR _10186_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13427__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13945_ _13944_/B _13946_/B _13944_/C _13944_/D VGND VGND VPWR VPWR _12992_/A sky130_fd_sc_hd__and4b_4
XFILLER_46_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ _13882_/CLK line[125] VGND VGND VPWR VPWR _13876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12827_ _12826_/Q _12852_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12774_/CLK line[126] VGND VGND VPWR VPWR _12759_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07160__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11709_ _11708_/Q _11732_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ _12688_/Q _12712_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_05230_ _05229_/Q _05257_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05161_ _05157_/CLK line[109] VGND VGND VPWR VPWR _05162_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09087__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05092_ _05091_/Q _05117_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[0\].VALID\[7\].TOBUF OVHB\[0\].VALID\[7\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_08920_ _08922_/CLK line[21] VGND VGND VPWR VPWR _08920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10026__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08851_ _08851_/A _08862_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12241__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07802_ _07788_/CLK line[22] VGND VGND VPWR VPWR _07802_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13915__A A[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04959__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05994_ _05993_/Q _06027_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_08782_ _08762_/CLK line[86] VGND VGND VPWR VPWR _08783_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07335__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07733_ _07732_/Q _07742_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_04945_ _04947_/CLK line[10] VGND VGND VPWR VPWR _04946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07664_ _07644_/CLK line[87] VGND VGND VPWR VPWR _07665_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09550__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09403_ _09402_/Q _09422_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06615_ _06615_/A _06622_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_07595_ _07595_/A _07602_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[29\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06546_ _06528_/CLK line[88] VGND VGND VPWR VPWR _06546_/Q sky130_fd_sc_hd__dfxtp_1
X_09334_ _09320_/CLK line[82] VGND VGND VPWR VPWR _09334_/Q sky130_fd_sc_hd__dfxtp_1
X_06477_ _06477_/A _06482_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_09265_ _09264_/Q _09282_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13800__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05428_ _05424_/CLK line[89] VGND VGND VPWR VPWR _05428_/Q sky130_fd_sc_hd__dfxtp_1
X_08216_ _08208_/CLK line[83] VGND VGND VPWR VPWR _08216_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VOBUF OVHB\[3\].V/Q OVHB\[3\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_09196_ _09200_/CLK line[19] VGND VGND VPWR VPWR _09197_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05359_ _05358_/Q _05362_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_08147_ _08147_/A _08162_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12416__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08078_ _08070_/CLK line[20] VGND VGND VPWR VPWR _08079_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07029_ _07029_/A _07042_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13097__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09725__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10040_ _10042_/CLK line[21] VGND VGND VPWR VPWR _10040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[31\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _11905_/CLK sky130_fd_sc_hd__clkbuf_4
X_11991_ _11990_/Q _12012_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11990__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ _13746_/CLK line[58] VGND VGND VPWR VPWR _13730_/Q sky130_fd_sc_hd__dfxtp_1
X_10942_ _10930_/CLK line[49] VGND VGND VPWR VPWR _10942_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09460__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13661_ _13660_/Q _13692_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_10873_ _10872_/Q _10892_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[9\].TOBUF OVHB\[31\].VALID\[9\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ _12638_/CLK line[59] VGND VGND VPWR VPWR _12613_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08076__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ _13598_/CLK line[123] VGND VGND VPWR VPWR _13592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[9\].VALID\[2\].TOBUF OVHB\[9\].VALID\[2\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ _12543_/A _12572_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12474_ _12490_/CLK line[124] VGND VGND VPWR VPWR _12474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11425_ _11424_/Q _11452_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11230__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _05150_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06324__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11356_ _11370_/CLK line[125] VGND VGND VPWR VPWR _11356_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06902__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ _10307_/A _10332_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_11287_ _11286_/Q _11312_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09635__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06621__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13026_ _12992_/A wr VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__and2_1
X_10238_ _10248_/CLK line[126] VGND VGND VPWR VPWR _10238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13157__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10169_ _10168_/Q _10192_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[27\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13928_ _13933_/B _13934_/B _13934_/C _13934_/D VGND VGND VPWR VPWR _09632_/A sky130_fd_sc_hd__nor4b_4
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13859_ _13845_/CLK line[103] VGND VGND VPWR VPWR _13860_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11405__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _11520_/CLK sky130_fd_sc_hd__clkbuf_4
X_06400_ _06408_/CLK line[21] VGND VGND VPWR VPWR _06400_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[10\].FF OVHB\[12\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[12\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07380_ _07380_/CLK line[85] VGND VGND VPWR VPWR _07381_/A sky130_fd_sc_hd__dfxtp_1
X_06331_ _06330_/Q _06342_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09050_ _09068_/CLK line[95] VGND VGND VPWR VPWR _09050_/Q sky130_fd_sc_hd__dfxtp_1
X_06262_ _06244_/CLK line[86] VGND VGND VPWR VPWR _06262_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08714__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08001_ _08001_/A _08022_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_05213_ _05212_/Q _05222_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06193_ _06192_/Q _06202_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[4\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11140__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05144_ _05122_/CLK line[87] VGND VGND VPWR VPWR _05145_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05075_ _05074_/Q _05082_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_09952_ _09978_/CLK line[123] VGND VGND VPWR VPWR _09952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[12\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08903_ _08902_/Q _08932_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_09883_ _09882_/Q _09912_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13067__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08834_ _08850_/CLK line[124] VGND VGND VPWR VPWR _08835_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07065__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08765_ _08765_/A _08792_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_05977_ _05977_/A _05992_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_07716_ _07724_/CLK line[125] VGND VGND VPWR VPWR _07717_/A sky130_fd_sc_hd__dfxtp_1
X_04928_ _04917_/Y _04918_/A2 A_h[12] _04927_/Y VGND VGND VPWR VPWR _04928_/X sky130_fd_sc_hd__a2bb2o_4
X_08696_ _08710_/CLK line[61] VGND VGND VPWR VPWR _08696_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07647_ _07646_/Q _07672_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11315__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[1\].FF OVHB\[21\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[21\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05313__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07578_ _07572_/CLK line[62] VGND VGND VPWR VPWR _07578_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[14\].TOBUF OVHB\[11\].VALID\[14\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_09317_ _09352_/A VGND VGND VPWR VPWR _09317_/Y sky130_fd_sc_hd__inv_2
X_06529_ _06528_/Q _06552_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13530__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _09256_/CLK line[48] VGND VGND VPWR VPWR _09248_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08624__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[27\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12146__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09179_ _09178_/Q _09212_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].CG clk OVHB\[22\].CGAND/X VGND VGND VPWR VPWR OVHB\[22\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_108_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11210_ _11216_/CLK line[58] VGND VGND VPWR VPWR _11210_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12190_ _12204_/CLK line[122] VGND VGND VPWR VPWR _12190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11141_ _11140_/Q _11172_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11072_ _11090_/CLK line[123] VGND VGND VPWR VPWR _11073_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10023_ _10023_/A _10052_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[7\].VALID\[7\].TOBUF OVHB\[7\].VALID\[7\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13705__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11974_ _11973_/Q _11977_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07703__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09190__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13713_ _13701_/CLK line[36] VGND VGND VPWR VPWR _13713_/Q sky130_fd_sc_hd__dfxtp_1
X_10925_ _10925_/CLK _10926_/X VGND VGND VPWR VPWR _10903_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_44_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[13\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _13643_/Q _13657_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_10856_ _11032_/A wr VGND VGND VPWR VPWR _10856_/X sky130_fd_sc_hd__and2_1
XANTENNA__05223__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13559_/CLK line[101] VGND VGND VPWR VPWR _13575_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ _13932_/X VGND VGND VPWR VPWR _10787_/Y sky130_fd_sc_hd__inv_2
XOVHB\[7\].VALID\[12\].FF OVHB\[7\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[7\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _12526_/A _12537_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12056__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12457_ _12449_/CLK line[102] VGND VGND VPWR VPWR _12457_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06054__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11408_ _11407_/Q _11417_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[27\]_A3 _13593_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12388_ _12388_/A _12397_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11895__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[0\].V OVHB\[0\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[0\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[0\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11339_ _11343_/CLK line[103] VGND VGND VPWR VPWR _11339_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06989__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[23\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09365__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05900_ _05902_/CLK line[63] VGND VGND VPWR VPWR _05900_/Q sky130_fd_sc_hd__dfxtp_1
X_13009_ _12999_/CLK line[98] VGND VGND VPWR VPWR _13009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10304__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06880_ _06892_/CLK line[127] VGND VGND VPWR VPWR _06880_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[14\].TOBUF OVHB\[31\].VALID\[14\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_05831_ _05830_/Q _05852_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_08550_ _08560_/CLK line[122] VGND VGND VPWR VPWR _08550_/Q sky130_fd_sc_hd__dfxtp_1
X_05762_ _05756_/CLK line[113] VGND VGND VPWR VPWR _05763_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07613__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07501_ _07500_/Q _07532_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08481_ _08481_/A _08512_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_05693_ _05693_/A _05712_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[14\].VALID\[2\].TOBUF OVHB\[14\].VALID\[2\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_07432_ _07446_/CLK line[123] VGND VGND VPWR VPWR _07432_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06229__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05711__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07363_ _07362_/Q _07392_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09102_ _09102_/A _09107_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_06314_ _06320_/CLK line[124] VGND VGND VPWR VPWR _06314_/Q sky130_fd_sc_hd__dfxtp_1
X_07294_ _07292_/CLK line[60] VGND VGND VPWR VPWR _07294_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[4\].FF OVHB\[18\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[18\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09033_ _09005_/CLK line[73] VGND VGND VPWR VPWR _09033_/Q sky130_fd_sc_hd__dfxtp_1
X_06245_ _06244_/Q _06272_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06176_ _06186_/CLK line[61] VGND VGND VPWR VPWR _06177_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05127_ _05126_/Q _05152_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09935_ _09925_/CLK line[101] VGND VGND VPWR VPWR _09935_/Q sky130_fd_sc_hd__dfxtp_1
X_05058_ _05058_/CLK line[62] VGND VGND VPWR VPWR _05058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09866_ _09865_/Q _09877_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08817_ _08823_/CLK line[102] VGND VGND VPWR VPWR _08817_/Q sky130_fd_sc_hd__dfxtp_1
X_09797_ _09793_/CLK line[38] VGND VGND VPWR VPWR _09798_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[3\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08748_ _08748_/A _08757_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08679_ _08663_/CLK line[39] VGND VGND VPWR VPWR _08680_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11045__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10709_/Q _10717_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06139__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05043__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11690_ _11690_/A _11697_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10641_ _10627_/CLK line[40] VGND VGND VPWR VPWR _10642_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05978__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13260__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ _13360_/A _13377_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08354__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10572_ _10572_/A _10577_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08932__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12311_ _12311_/CLK line[35] VGND VGND VPWR VPWR _12311_/Q sky130_fd_sc_hd__dfxtp_1
X_13291_ _13285_/CLK line[99] VGND VGND VPWR VPWR _13291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08651__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12242_ _12241_/Q _12257_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[1\].TOBUF OVHB\[20\].VALID\[1\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_123_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12173_ _12177_/CLK line[100] VGND VGND VPWR VPWR _12173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[16\].VALID\[6\].FF OVHB\[16\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[16\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11124_ _11123_/Q _11137_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06602__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11055_ _11063_/CLK line[101] VGND VGND VPWR VPWR _11056_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09913__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05218__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10006_ _10005_/Q _10017_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13435__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08529__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11957_ _11945_/CLK line[1] VGND VGND VPWR VPWR _11957_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08826__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10908_ _10907_/Q _10927_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_11888_ _11887_/Q _11907_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13627_ _13631_/CLK line[11] VGND VGND VPWR VPWR _13627_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10794__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10839_ _10843_/CLK line[2] VGND VGND VPWR VPWR _10840_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13170__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05888__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13558_ _13557_/Q _13587_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_12509_ _12523_/CLK line[12] VGND VGND VPWR VPWR _12509_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].INV _13967_/X VGND VGND VPWR VPWR OVHB\[22\].INV/Y sky130_fd_sc_hd__inv_2
X_13489_ _13497_/CLK line[76] VGND VGND VPWR VPWR _13489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06030_ _06050_/CLK line[122] VGND VGND VPWR VPWR _06031_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09095__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07981_ _07981_/CLK line[104] VGND VGND VPWR VPWR _07982_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[12\].VALID\[7\].TOBUF OVHB\[12\].VALID\[7\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09720_ _09719_/Q _09737_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10034__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06932_ _06932_/A _06937_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10612__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05128__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09651_ _09659_/CLK line[99] VGND VGND VPWR VPWR _09652_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10969__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06863_ _06839_/CLK line[105] VGND VGND VPWR VPWR _06863_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10331__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[11\].TOBUF OVHB\[5\].VALID\[11\].FF/Q OVHB\[5\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13345__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08602_ _08601_/Q _08617_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_05814_ _05813_/Q _05817_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04967__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09582_ _09581_/Q _09597_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[8\].FF OVHB\[14\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[14\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07343__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06794_ _06793_/Q _06797_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[10\].FF OVHB\[3\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[3\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08533_ _08541_/CLK line[100] VGND VGND VPWR VPWR _08533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05745_ _05745_/CLK _05746_/X VGND VGND VPWR VPWR _05739_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _08464_/A _08477_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05676_ _13909_/X wr VGND VGND VPWR VPWR _05676_/X sky130_fd_sc_hd__and2_1
X_07415_ _07393_/CLK line[101] VGND VGND VPWR VPWR _07415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _08383_/CLK line[37] VGND VGND VPWR VPWR _08395_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07346_ _07345_/Q _07357_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10209__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07277_ _07267_/CLK line[38] VGND VGND VPWR VPWR _07277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09016_ _09016_/A _09037_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_06228_ _06227_/Q _06237_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08902__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06272__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10506__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06159_ _06147_/CLK line[39] VGND VGND VPWR VPWR _06159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12424__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07518__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09918_ _09918_/A _09947_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09733__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09849_ _09849_/CLK line[76] VGND VGND VPWR VPWR _09849_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[9\]_A3 _06864_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12860_ _12859_/Q _12887_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07253__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11811_ _11823_/CLK line[77] VGND VGND VPWR VPWR _11811_/Q sky130_fd_sc_hd__dfxtp_1
X_12791_ _12803_/CLK line[13] VGND VGND VPWR VPWR _12791_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[17\]_A2 _06533_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11742_ _11741_/Q _11767_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06447__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11691_/CLK line[14] VGND VGND VPWR VPWR _11673_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06166__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13552_/A VGND VGND VPWR VPWR _13412_/Y sky130_fd_sc_hd__inv_2
X_10624_ _10623_/Q _10647_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08084__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[13\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13343_ _13347_/CLK line[0] VGND VGND VPWR VPWR _13343_/Q sky130_fd_sc_hd__dfxtp_1
X_10555_ _10571_/CLK line[15] VGND VGND VPWR VPWR _10555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09908__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13274_ _13273_/Q _13307_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_10486_ _10485_/Q _10507_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12334__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12225_ _12227_/CLK line[10] VGND VGND VPWR VPWR _12225_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07428__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06332__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12156_ _12156_/A _12187_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11107_ _11111_/CLK line[11] VGND VGND VPWR VPWR _11108_/A sky130_fd_sc_hd__dfxtp_1
X_12087_ _12109_/CLK line[75] VGND VGND VPWR VPWR _12087_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09643__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11038_ _11037_/Q _11067_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[10\].FF OVHB\[17\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[17\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08259__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07741__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12989_ _12988_/Q _12992_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[13\].TOBUF OVHB\[28\].VALID\[13\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_05530_ _05530_/A _05537_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05461_ _05445_/CLK line[104] VGND VGND VPWR VPWR _05462_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12509__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11413__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07200_ _07199_/Q _07217_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05392_ _05391_/Q _05397_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_08180_ _08179_/Q _08197_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06507__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07131_ _07117_/CLK line[99] VGND VGND VPWR VPWR _07132_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09818__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07062_ _07062_/A _07077_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_06013_ _06023_/CLK line[100] VGND VGND VPWR VPWR _06013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06242__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[1\].TOBUF OVHB\[27\].VALID\[1\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07964_ _07963_/Q _07987_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[12\].TOBUF OVHB\[21\].VALID\[12\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_68_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09703_ _09721_/CLK line[0] VGND VGND VPWR VPWR _09703_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10699__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06915_ _06923_/CLK line[15] VGND VGND VPWR VPWR _06916_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07895_ _07905_/CLK line[79] VGND VGND VPWR VPWR _07895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13075__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09634_ _09633_/Q _09667_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_06846_ _06846_/A _06867_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08169__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07073__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10996__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09565_ _09577_/CLK line[74] VGND VGND VPWR VPWR _09565_/Q sky130_fd_sc_hd__dfxtp_1
X_06777_ _06775_/CLK line[65] VGND VGND VPWR VPWR _06778_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[1\].FF OVHB\[7\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[7\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08516_ _08515_/Q _08547_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05728_ _05727_/Q _05747_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _09495_/Q _09527_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _08473_/CLK line[75] VGND VGND VPWR VPWR _08447_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[26\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05659_ _05671_/CLK line[66] VGND VGND VPWR VPWR _05659_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11323__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06417__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _08377_/Q _08407_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05321__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07329_ _07327_/CLK line[76] VGND VGND VPWR VPWR _07330_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10340_ _10339_/Q _10367_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08632__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[19\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10271_ _10277_/CLK line[13] VGND VGND VPWR VPWR _10271_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07248__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12010_ _12010_/CLK _12011_/X VGND VGND VPWR VPWR _12002_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04938__B2 _04938_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13961_ _13958_/X _13964_/B _13960_/X _13966_/D VGND VGND VPWR VPWR _13961_/Y sky130_fd_sc_hd__nor4b_4
XFILLER_98_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[19\].VALID\[7\].TOBUF OVHB\[19\].VALID\[7\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12912_ _12902_/CLK line[54] VGND VGND VPWR VPWR _12912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13892_ _13882_/CLK line[118] VGND VGND VPWR VPWR _13893_/A sky130_fd_sc_hd__dfxtp_1
X_12843_ _12842_/Q _12852_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13713__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08807__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12774_ _12774_/CLK line[119] VGND VGND VPWR VPWR _12774_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05081__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11725_ _11725_/A _11732_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11656_ _11636_/CLK line[120] VGND VGND VPWR VPWR _11657_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05231__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[7\].INV _13990_/X VGND VGND VPWR VPWR OVHB\[7\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[3\].FF OVHB\[5\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[5\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10607_ _10606_/Q _10612_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11586_/Q _11592_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_13326_ _13308_/CLK line[115] VGND VGND VPWR VPWR _13326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10538_ _10520_/CLK line[121] VGND VGND VPWR VPWR _10538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12064__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13257_ _13256_/Q _13272_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12642__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10469_ _10469_/A _10472_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].V OVHB\[27\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[27\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07158__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12208_ _12204_/CLK line[116] VGND VGND VPWR VPWR _12208_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12999__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13188_ _13194_/CLK line[52] VGND VGND VPWR VPWR _13188_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12361__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06997__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12139_ _12138_/Q _12152_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09373__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05256__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04961_ _04947_/CLK line[3] VGND VGND VPWR VPWR _04961_/Q sky130_fd_sc_hd__dfxtp_1
X_06700_ _06700_/A _06727_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10312__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07680_ _07680_/A _07707_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05406__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06631_ _06633_/CLK line[13] VGND VGND VPWR VPWR _06632_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13623__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09350_ _09350_/CLK _09351_/X VGND VGND VPWR VPWR _09320_/CLK sky130_fd_sc_hd__dlclkp_1
X_06562_ _06561_/Q _06587_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[3\].TOBUF OVHB\[0\].VALID\[3\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__07621__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08301_ _13940_/X wr VGND VGND VPWR VPWR _08301_/X sky130_fd_sc_hd__and2_1
X_05513_ _05519_/CLK line[14] VGND VGND VPWR VPWR _05513_/Q sky130_fd_sc_hd__dfxtp_1
X_09281_ _09352_/A wr VGND VGND VPWR VPWR _09281_/X sky130_fd_sc_hd__and2_1
XANTENNA__12239__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06493_ _06489_/CLK line[78] VGND VGND VPWR VPWR _06493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12817__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[6\].TOBUF OVHB\[25\].VALID\[6\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_08232_ _13940_/X VGND VGND VPWR VPWR _08232_/Y sky130_fd_sc_hd__inv_2
X_05444_ _05443_/Q _05467_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12536__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08163_ _08175_/CLK line[64] VGND VGND VPWR VPWR _08163_/Q sky130_fd_sc_hd__dfxtp_1
X_05375_ _05391_/CLK line[79] VGND VGND VPWR VPWR _05375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09548__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07114_ _07113_/Q _07147_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04980__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08094_ _08093_/Q _08127_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_07045_ _07043_/CLK line[74] VGND VGND VPWR VPWR _07046_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].V OVHB\[18\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[18\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[3\].VALID\[5\].FF OVHB\[3\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[3\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12702__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08996_ _08972_/CLK line[56] VGND VGND VPWR VPWR _08996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09283__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07947_ _07947_/A _07952_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07878_ _07854_/CLK line[57] VGND VGND VPWR VPWR _07879_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08477__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09617_ _09616_/Q _09632_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06829_ _06829_/A _06832_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08196__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09548_ _09554_/CLK line[52] VGND VGND VPWR VPWR _09549_/A sky130_fd_sc_hd__dfxtp_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XMUX.MUX\[31\] _10871_/Z _13461_/Z _11851_/Z _13601_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[31] sky130_fd_sc_hd__mux4_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _09478_/Q _09492_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ _11500_/CLK line[53] VGND VGND VPWR VPWR _11510_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06147__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12490_/CLK line[117] VGND VGND VPWR VPWR _12491_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11988__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _11440_/Q _11452_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05986__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09458__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08362__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11372_ _11370_/CLK line[118] VGND VGND VPWR VPWR _11372_/Q sky130_fd_sc_hd__dfxtp_1
X_13111_ _13110_/Q _13132_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_10323_ _10322_/Q _10332_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[31\].VALID\[5\].TOBUF OVHB\[31\].VALID\[5\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_13042_ _13050_/CLK line[113] VGND VGND VPWR VPWR _13042_/Q sky130_fd_sc_hd__dfxtp_1
X_10254_ _10248_/CLK line[119] VGND VGND VPWR VPWR _10255_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12612__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10185_ _10184_/Q _10192_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06610__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09771__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11228__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13944_ _13946_/B _13944_/B _13944_/C _13944_/D VGND VGND VPWR VPWR _12712_/A sky130_fd_sc_hd__and4b_4
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09921__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[7\].FF OVHB\[1\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[1\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13875_ _13875_/A _13902_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13443__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12826_ _12820_/CLK line[29] VGND VGND VPWR VPWR _12826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08537__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12757_ _12756_/Q _12782_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11706_/CLK line[30] VGND VGND VPWR VPWR _11708_/Q sky130_fd_sc_hd__dfxtp_1
X_12688_ _12708_/CLK line[94] VGND VGND VPWR VPWR _12688_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11639_ _11639_/A _11662_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[16\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10157__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05896__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05160_ _05159_/Q _05187_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08272__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09946__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13309_ _13309_/A _13342_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
X_05091_ _05093_/CLK line[77] VGND VGND VPWR VPWR _05091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13618__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08850_ _08850_/CLK line[117] VGND VGND VPWR VPWR _08851_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[10\].FF OVHB\[8\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[8\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07801_ _07800_/Q _07812_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06520__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08781_ _08780_/Q _08792_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_05993_ _06023_/CLK line[96] VGND VGND VPWR VPWR _05993_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11138__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10042__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07732_ _07724_/CLK line[118] VGND VGND VPWR VPWR _07732_/Q sky130_fd_sc_hd__dfxtp_1
X_04944_ _04943_/Q _04977_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05136__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10977__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07663_ _07663_/A _07672_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[11\].TOBUF OVHB\[18\].VALID\[11\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13353__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09402_ _09414_/CLK line[113] VGND VGND VPWR VPWR _09402_/Q sky130_fd_sc_hd__dfxtp_1
X_06614_ _06596_/CLK line[119] VGND VGND VPWR VPWR _06615_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[22\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08447__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07594_ _07572_/CLK line[55] VGND VGND VPWR VPWR _07595_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07351__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09333_ _09333_/A _09352_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_06545_ _06544_/Q _06552_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11451__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09264_ _09256_/CLK line[50] VGND VGND VPWR VPWR _09264_/Q sky130_fd_sc_hd__dfxtp_1
X_06476_ _06464_/CLK line[56] VGND VGND VPWR VPWR _06477_/A sky130_fd_sc_hd__dfxtp_1
X_08215_ _08215_/A _08232_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_05427_ _05427_/A _05432_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09195_ _09195_/A _09212_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11601__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09278__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08146_ _08134_/CLK line[51] VGND VGND VPWR VPWR _08147_/A sky130_fd_sc_hd__dfxtp_1
X_05358_ _05332_/CLK line[57] VGND VGND VPWR VPWR _05358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10217__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08077_ _08076_/Q _08092_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_05289_ _05289_/A _05292_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07028_ _07030_/CLK line[52] VGND VGND VPWR VPWR _07029_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08910__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13528__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[10\].TOBUF OVHB\[11\].VALID\[10\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07526__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[2\].FF OVHB\[28\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[28\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08979_ _08978_/Q _09002_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11626__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].CGAND _12992_/A wr VGND VGND VPWR VPWR OVHB\[6\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_57_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11990_ _12002_/CLK line[31] VGND VGND VPWR VPWR _11990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10941_ _10940_/Q _10962_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13660_ _13682_/CLK line[26] VGND VGND VPWR VPWR _13660_/Q sky130_fd_sc_hd__dfxtp_1
X_10872_ _10872_/CLK line[17] VGND VGND VPWR VPWR _10872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07261__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ _12610_/Q _12642_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ _13590_/Q _13622_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _12560_/CLK line[27] VGND VGND VPWR VPWR _12543_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[3\].TOBUF OVHB\[7\].VALID\[3\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12473_ _12472_/Q _12502_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09188__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11424_ _11440_/CLK line[28] VGND VGND VPWR VPWR _11424_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10127__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11355_ _11354_/Q _11382_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07286__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10306_ _10314_/CLK line[29] VGND VGND VPWR VPWR _10307_/A sky130_fd_sc_hd__dfxtp_1
X_11286_ _11302_/CLK line[93] VGND VGND VPWR VPWR _11286_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12342__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13025_ _13025_/CLK _13026_/X VGND VGND VPWR VPWR _12999_/CLK sky130_fd_sc_hd__dlclkp_1
X_10237_ _10236_/Q _10262_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07436__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10168_ _10188_/CLK line[94] VGND VGND VPWR VPWR _10168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10099_ _10098_/Q _10122_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09651__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13927_ A[6] VGND VGND VPWR VPWR _13934_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_90_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ _13857_/Q _13867_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[26\].VALID\[4\].FF OVHB\[26\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[26\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12809_ _12803_/CLK line[7] VGND VGND VPWR VPWR _12810_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13789_ _13763_/CLK line[71] VGND VGND VPWR VPWR _13789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[28\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06330_ _06320_/CLK line[117] VGND VGND VPWR VPWR _06330_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12517__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06261_ _06260_/Q _06272_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _10890_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[31\].VALID\[10\].TOBUF OVHB\[31\].VALID\[10\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_08000_ _08000_/CLK line[127] VGND VGND VPWR VPWR _08001_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[2\].CGAND_A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05212_ _05214_/CLK line[118] VGND VGND VPWR VPWR _05212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06192_ _06186_/CLK line[54] VGND VGND VPWR VPWR _06192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[19\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _08020_/CLK sky130_fd_sc_hd__clkbuf_4
X_05143_ _05142_/Q _05152_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09826__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05074_ _05058_/CLK line[55] VGND VGND VPWR VPWR _05074_/Q sky130_fd_sc_hd__dfxtp_1
X_09951_ _09951_/A _09982_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_MUX.MUX\[12\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[14\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08902_ _08922_/CLK line[27] VGND VGND VPWR VPWR _08902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13926__A A[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09882_ _09908_/CLK line[91] VGND VGND VPWR VPWR _09882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08833_ _08832_/Q _08862_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06250__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08764_ _08762_/CLK line[92] VGND VGND VPWR VPWR _08765_/A sky130_fd_sc_hd__dfxtp_1
X_05976_ _05984_/CLK line[83] VGND VGND VPWR VPWR _05977_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[7\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07715_ _07714_/Q _07742_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_04927_ _04927_/A VGND VGND VPWR VPWR _04927_/Y sky130_fd_sc_hd__inv_2
X_08695_ _08694_/Q _08722_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13083__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08177__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07646_ _07644_/CLK line[93] VGND VGND VPWR VPWR _07646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07577_ _07576_/Q _07602_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09316_ _09352_/A wr VGND VGND VPWR VPWR _09316_/X sky130_fd_sc_hd__and2_1
X_06528_ _06528_/CLK line[94] VGND VGND VPWR VPWR _06528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[7\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09247_ _09352_/A VGND VGND VPWR VPWR _09247_/Y sky130_fd_sc_hd__inv_2
X_06459_ _06458_/Q _06482_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11331__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[6\].FF OVHB\[24\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[24\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06425__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09178_ _09200_/CLK line[16] VGND VGND VPWR VPWR _09178_/Q sky130_fd_sc_hd__dfxtp_1
X_08129_ _08128_/Q _08162_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_11140_ _11148_/CLK line[26] VGND VGND VPWR VPWR _11140_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08640__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13258__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11071_ _11070_/Q _11102_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[18\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _07635_/CLK sky130_fd_sc_hd__clkbuf_4
X_10022_ _10042_/CLK line[27] VGND VGND VPWR VPWR _10023_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[8\].TOBUF OVHB\[5\].VALID\[8\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_11973_ _11945_/CLK line[9] VGND VGND VPWR VPWR _11973_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11506__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13712_ _13711_/Q _13727_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_10924_ _10924_/A _10927_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13643_ _13631_/CLK line[4] VGND VGND VPWR VPWR _13643_/Q sky130_fd_sc_hd__dfxtp_1
X_10855_ _10855_/CLK _10856_/X VGND VGND VPWR VPWR _10843_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12187__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13721__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08815__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13574_ _13573_/Q _13587_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _13932_/X wr VGND VGND VPWR VPWR _10786_/X sky130_fd_sc_hd__and2_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _12523_/CLK line[5] VGND VGND VPWR VPWR _12526_/A sky130_fd_sc_hd__dfxtp_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12456_ _12455_/Q _12467_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_11407_ _11395_/CLK line[6] VGND VGND VPWR VPWR _11407_/Q sky130_fd_sc_hd__dfxtp_1
X_12387_ _12387_/CLK line[70] VGND VGND VPWR VPWR _12388_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11338_ _11337_/Q _11347_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08550__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13168__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12072__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11269_ _11251_/CLK line[71] VGND VGND VPWR VPWR _11269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07166__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[8\].FF OVHB\[22\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[22\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13008_ _13007_/Q _13027_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[13\].FF OVHB\[30\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[30\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05830_ _05836_/CLK line[31] VGND VGND VPWR VPWR _05830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09381__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _07250_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_48_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05761_ _05761_/A _05782_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13481__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07500_ _07518_/CLK line[26] VGND VGND VPWR VPWR _07500_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10320__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08480_ _08480_/CLK line[90] VGND VGND VPWR VPWR _08481_/A sky130_fd_sc_hd__dfxtp_1
X_05692_ _05708_/CLK line[81] VGND VGND VPWR VPWR _05693_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05414__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07431_ _07430_/Q _07462_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13631__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[3\].TOBUF OVHB\[12\].VALID\[3\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__08725__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07362_ _07380_/CLK line[91] VGND VGND VPWR VPWR _07362_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05711__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09101_ _09085_/CLK line[104] VGND VGND VPWR VPWR _09102_/A sky130_fd_sc_hd__dfxtp_1
X_06313_ _06312_/Q _06342_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12247__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07293_ _07292_/Q _07322_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ _09031_/Q _09037_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_06244_ _06244_/CLK line[92] VGND VGND VPWR VPWR _06244_/Q sky130_fd_sc_hd__dfxtp_1
X_06175_ _06174_/Q _06202_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09556__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05126_ _05122_/CLK line[93] VGND VGND VPWR VPWR _05126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13656__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09934_ _09933_/Q _09947_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_05057_ _05056_/Q _05082_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09865_ _09849_/CLK line[69] VGND VGND VPWR VPWR _09865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13806__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08816_ _08815_/Q _08827_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_09796_ _09795_/Q _09807_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09291__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07804__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[12\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08747_ _08749_/CLK line[70] VGND VGND VPWR VPWR _08748_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05959_ _05958_/Q _05992_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10230__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08678_ _08677_/Q _08687_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DECH.DEC0.AND2_A_N A_h[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07633_/CLK line[71] VGND VGND VPWR VPWR _07629_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10640_/A _10647_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12157__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10571_ _10571_/CLK line[8] VGND VGND VPWR VPWR _10572_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11061__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12310_ _12309_/Q _12327_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06155__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13290_ _13289_/Q _13307_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11996__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12241_ _12227_/CLK line[3] VGND VGND VPWR VPWR _12241_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[5\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09466__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12172_ _12171_/Q _12187_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_11123_ _11111_/CLK line[4] VGND VGND VPWR VPWR _11123_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10405__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11054_ _11053_/Q _11067_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10005_ _10011_/CLK line[5] VGND VGND VPWR VPWR _10005_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12620__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07714__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[8\].VALID\[13\].TOBUF OVHB\[8\].VALID\[13\].FF/Q OVHB\[8\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_17_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11236__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11956_ _11955_/Q _11977_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_10907_ _10903_/CLK line[33] VGND VGND VPWR VPWR _10907_/Q sky130_fd_sc_hd__dfxtp_1
X_11887_ _11901_/CLK line[97] VGND VGND VPWR VPWR _11887_/Q sky130_fd_sc_hd__dfxtp_1
XMUX.MUX\[6\] _09448_/Z _05038_/Z _13508_/Z _13578_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[6] sky130_fd_sc_hd__mux4_1
X_13626_ _13625_/Q _13657_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_10838_ _10837_/Q _10857_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_10769_ _10783_/CLK line[98] VGND VGND VPWR VPWR _10770_/A sky130_fd_sc_hd__dfxtp_1
X_13557_ _13559_/CLK line[107] VGND VGND VPWR VPWR _13557_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06065__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12508_ _12507_/Q _12537_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
X_13488_ _13487_/Q _13517_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_12439_ _12449_/CLK line[108] VGND VGND VPWR VPWR _12439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08280__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[1\].VALID\[12\].TOBUF OVHB\[1\].VALID\[12\].FF/Q OVHB\[1\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_07980_ _07979_/Q _07987_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[14\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06931_ _06923_/CLK line[8] VGND VGND VPWR VPWR _06932_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[8\].TOBUF OVHB\[10\].VALID\[8\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_80_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09650_ _09650_/A _09667_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
X_06862_ _06862_/A _06867_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08601_ _08609_/CLK line[3] VGND VGND VPWR VPWR _08601_/Q sky130_fd_sc_hd__dfxtp_1
X_05813_ _05799_/CLK line[9] VGND VGND VPWR VPWR _05813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09581_ _09577_/CLK line[67] VGND VGND VPWR VPWR _09581_/Q sky130_fd_sc_hd__dfxtp_1
X_06793_ _06775_/CLK line[73] VGND VGND VPWR VPWR _06793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11146__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08532_ _08532_/A _08547_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_05744_ _05744_/A _05747_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].CG clk OVHB\[12\].CGAND/X VGND VGND VPWR VPWR OVHB\[12\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05144__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ _08473_/CLK line[68] VGND VGND VPWR VPWR _08464_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10985__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05675_ _05675_/CLK _05676_/X VGND VGND VPWR VPWR _05671_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13361__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07414_ _07413_/Q _07427_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08455__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ _08393_/Q _08407_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07345_ _07327_/CLK line[69] VGND VGND VPWR VPWR _07345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07276_ _07276_/A _07287_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09015_ _09005_/CLK line[79] VGND VGND VPWR VPWR _09016_/A sky130_fd_sc_hd__dfxtp_1
X_06227_ _06223_/CLK line[70] VGND VGND VPWR VPWR _06227_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06703__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06158_ _06158_/A _06167_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_05109_ _05093_/CLK line[71] VGND VGND VPWR VPWR _05109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06089_ _06077_/CLK line[7] VGND VGND VPWR VPWR _06090_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05319__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09917_ _09925_/CLK line[107] VGND VGND VPWR VPWR _09918_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13536__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[26\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09848_ _09847_/Q _09877_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09779_ _09793_/CLK line[44] VGND VGND VPWR VPWR _09780_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[25\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11810_ _11809_/Q _11837_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_12790_ _12789_/Q _12817_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05054__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[17\]_A3 _05203_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11741_ _11757_/CLK line[45] VGND VGND VPWR VPWR _11741_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10895__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11671_/Q _11697_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[14\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _10627_/CLK line[46] VGND VGND VPWR VPWR _10623_/Q sky130_fd_sc_hd__dfxtp_1
X_13411_ _13552_/A wr VGND VGND VPWR VPWR _13411_/X sky130_fd_sc_hd__and2_1
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _13272_/A VGND VGND VPWR VPWR _13342_/Y sky130_fd_sc_hd__inv_2
XOVHB\[19\].VALID\[3\].TOBUF OVHB\[19\].VALID\[3\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_10554_ _10553_/Q _10577_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_13273_ _13285_/CLK line[96] VGND VGND VPWR VPWR _13273_/Q sky130_fd_sc_hd__dfxtp_1
X_10485_ _10473_/CLK line[111] VGND VGND VPWR VPWR _10485_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09196__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12224_ _12223_/Q _12257_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[27\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _12177_/CLK line[106] VGND VGND VPWR VPWR _12156_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10135__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05229__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11106_ _11105_/Q _11137_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[24\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12086_ _12085_/Q _12117_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[24\].VALID\[14\].TOBUF OVHB\[24\].VALID\[14\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__12350__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11037_ _11063_/CLK line[107] VGND VGND VPWR VPWR _11037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07444__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07741__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12988_ _12962_/CLK line[89] VGND VGND VPWR VPWR _12988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[7\].CG clk OVHB\[7\].CGAND/X VGND VGND VPWR VPWR OVHB\[7\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_11939_ _11938_/Q _11942_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_05460_ _05460_/A _05467_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13609_ _13608_/Q _13622_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05391_ _05391_/CLK line[72] VGND VGND VPWR VPWR _05391_/Q sky130_fd_sc_hd__dfxtp_1
X_07130_ _07129_/Q _07147_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12525__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07061_ _07043_/CLK line[67] VGND VGND VPWR VPWR _07062_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07619__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06012_ _06011_/Q _06027_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09834__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07963_ _07981_/CLK line[110] VGND VGND VPWR VPWR _07963_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[2\].TOBUF OVHB\[25\].VALID\[2\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[8\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _13550_/CLK sky130_fd_sc_hd__clkbuf_4
X_06914_ _06913_/Q _06937_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_09702_ _09632_/A VGND VGND VPWR VPWR _09702_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12260__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__04978__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07894_ _07893_/Q _07917_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09633_ _09659_/CLK line[96] VGND VGND VPWR VPWR _09633_/Q sky130_fd_sc_hd__dfxtp_1
X_06845_ _06839_/CLK line[111] VGND VGND VPWR VPWR _06846_/A sky130_fd_sc_hd__dfxtp_1
X_09564_ _09563_/Q _09597_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_06776_ _06776_/A _06797_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08515_ _08541_/CLK line[106] VGND VGND VPWR VPWR _08515_/Q sky130_fd_sc_hd__dfxtp_1
X_05727_ _05739_/CLK line[97] VGND VGND VPWR VPWR _05727_/Q sky130_fd_sc_hd__dfxtp_1
X_09495_ _09507_/CLK line[42] VGND VGND VPWR VPWR _09495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13091__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08185__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08446_ _08445_/Q _08477_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05658_ _05658_/A _05677_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ _08383_/CLK line[43] VGND VGND VPWR VPWR _08377_/Q sky130_fd_sc_hd__dfxtp_1
X_05589_ _05575_/CLK line[34] VGND VGND VPWR VPWR _05589_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07328_ _07328_/A _07357_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12435__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07259_ _07267_/CLK line[44] VGND VGND VPWR VPWR _07259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06433__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10270_ _10269_/Q _10297_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09744__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13266__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13960_ A_h[6] VGND VGND VPWR VPWR _13960_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12911_ _12910_/Q _12922_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[8\].TOBUF OVHB\[17\].VALID\[8\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_13891_ _13890_/Q _13902_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].INV _13966_/X VGND VGND VPWR VPWR OVHB\[21\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_46_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12842_ _12820_/CLK line[22] VGND VGND VPWR VPWR _12842_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _13165_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13983__D_N _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05362__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[24\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12773_ _12772_/Q _12782_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[1\].TOBUF OVHB\[31\].VALID\[1\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11514__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08095__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05081__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06608__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11724_ _11706_/CLK line[23] VGND VGND VPWR VPWR _11725_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[30\]_A0 _09469_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11662_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09919__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08823__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10606_ _10594_/CLK line[24] VGND VGND VPWR VPWR _10606_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11588_/CLK line[88] VGND VGND VPWR VPWR _11586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13325_ _13324_/Q _13342_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_10537_ _10537_/A _10542_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06343__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10468_ _10466_/CLK line[89] VGND VGND VPWR VPWR _10469_/A sky130_fd_sc_hd__dfxtp_1
X_13256_ _13254_/CLK line[83] VGND VGND VPWR VPWR _13256_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[8\].FF OVHB\[8\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[8\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12207_ _12207_/A _12222_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_13187_ _13187_/A _13202_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10399_ _10398_/Q _10402_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05537__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _12130_/CLK line[84] VGND VGND VPWR VPWR _12138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13176__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[27\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _10505_/CLK sky130_fd_sc_hd__clkbuf_4
X_12069_ _12068_/Q _12082_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05256__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04960_ _04960_/A _04977_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07174__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06630_ _06629_/Q _06657_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06561_ _06565_/CLK line[109] VGND VGND VPWR VPWR _06561_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11424__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08300_ _08300_/CLK _08301_/X VGND VGND VPWR VPWR _08282_/CLK sky130_fd_sc_hd__dlclkp_1
X_05512_ _05511_/Q _05537_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06518__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09280_ _09280_/CLK _09281_/X VGND VGND VPWR VPWR _09256_/CLK sky130_fd_sc_hd__dlclkp_1
X_06492_ _06492_/A _06517_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05422__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08231_ _13940_/X wr VGND VGND VPWR VPWR _08231_/X sky130_fd_sc_hd__and2_1
X_05443_ _05445_/CLK line[110] VGND VGND VPWR VPWR _05443_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[7\].TOBUF OVHB\[23\].VALID\[7\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_127_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08162_ _13940_/X VGND VGND VPWR VPWR _08162_/Y sky130_fd_sc_hd__inv_2
XANTENNA_MUX.MUX\[7\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08733__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05374_ _05374_/A _05397_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_07113_ _07117_/CLK line[96] VGND VGND VPWR VPWR _07113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08093_ _08113_/CLK line[32] VGND VGND VPWR VPWR _08093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07349__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07044_ _07043_/Q _07077_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06831__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08995_ _08995_/A _09002_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10503__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07946_ _07946_/CLK line[88] VGND VGND VPWR VPWR _07947_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07084__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07877_ _07876_/Q _07882_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13814__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09616_ _09626_/CLK line[83] VGND VGND VPWR VPWR _09616_/Q sky130_fd_sc_hd__dfxtp_1
X_06828_ _06802_/CLK line[89] VGND VGND VPWR VPWR _06829_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[26\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _10120_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08908__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06759_ _06758_/Q _06762_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_09547_ _09546_/Q _09562_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05332__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09478_ _09482_/CLK line[20] VGND VGND VPWR VPWR _09478_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[24\] _10887_/Z _13477_/Z _13547_/Z _12777_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[24] sky130_fd_sc_hd__mux4_1
X_08429_ _08428_/Q _08442_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _11440_/CLK line[21] VGND VGND VPWR VPWR _11440_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[2\].CGAND _11311_/A wr VGND VGND VPWR VPWR OVHB\[2\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA_OVHB\[23\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12165__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11371_ _11371_/A _11382_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07259__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06163__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13110_ _13120_/CLK line[31] VGND VGND VPWR VPWR _13110_/Q sky130_fd_sc_hd__dfxtp_1
X_10322_ _10314_/CLK line[22] VGND VGND VPWR VPWR _10322_/Q sky130_fd_sc_hd__dfxtp_1
X_13041_ _13041_/A _13062_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_10253_ _10252_/Q _10262_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09474__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[16\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10184_ _10188_/CLK line[87] VGND VGND VPWR VPWR _10184_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[0\].FF OVHB\[17\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[17\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10413__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09771__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05507__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13943_ _13944_/B _13946_/B _13944_/C _13944_/D VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__and4bb_4
XFILLER_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13874_ _13882_/CLK line[124] VGND VGND VPWR VPWR _13875_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07722__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12825_ _12824_/Q _12852_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06338__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12774_/CLK line[125] VGND VGND VPWR VPWR _12756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[25\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _09735_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11706_/Q _11732_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12686_/Q _12712_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09649__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[15\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _06865_/CLK sky130_fd_sc_hd__clkbuf_4
X_11638_ _11636_/CLK line[126] VGND VGND VPWR VPWR _11639_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[22\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09946__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11569_ _11568_/Q _11592_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06073__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13308_ _13308_/CLK line[112] VGND VGND VPWR VPWR _13309_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05090_ _05090_/A _05117_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12803__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13239_ _13239_/A _13272_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[12\].TOBUF OVHB\[14\].VALID\[12\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_07800_ _07788_/CLK line[21] VGND VGND VPWR VPWR _07800_/Q sky130_fd_sc_hd__dfxtp_1
X_08780_ _08762_/CLK line[85] VGND VGND VPWR VPWR _08780_/Q sky130_fd_sc_hd__dfxtp_1
X_05992_ _13910_/X VGND VGND VPWR VPWR _05992_/Y sky130_fd_sc_hd__inv_2
X_07731_ _07730_/Q _07742_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_04943_ _04947_/CLK line[0] VGND VGND VPWR VPWR _04943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07662_ _07644_/CLK line[86] VGND VGND VPWR VPWR _07663_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[2\].FF OVHB\[15\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[15\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06613_ _06612_/Q _06622_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_09401_ _09400_/Q _09422_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07593_ _07592_/Q _07602_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11154__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11732__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06544_ _06528_/CLK line[87] VGND VGND VPWR VPWR _06544_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06248__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09332_ _09320_/CLK line[81] VGND VGND VPWR VPWR _09333_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[31\].VALID\[11\].FF OVHB\[31\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[31\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09263_ _09262_/Q _09282_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10993__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11451__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06475_ _06475_/A _06482_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08214_ _08208_/CLK line[82] VGND VGND VPWR VPWR _08215_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08463__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05426_ _05424_/CLK line[88] VGND VGND VPWR VPWR _05427_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ _09200_/CLK line[18] VGND VGND VPWR VPWR _09195_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08145_ _08144_/Q _08162_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_05357_ _05357_/A _05362_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_08076_ _08070_/CLK line[19] VGND VGND VPWR VPWR _08076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05288_ _05278_/CLK line[25] VGND VGND VPWR VPWR _05289_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[14\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _06480_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07027_ _07026_/Q _07042_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12713__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06711__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11329__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11907__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08978_ _08972_/CLK line[62] VGND VGND VPWR VPWR _08978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07392__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].INV _13989_/X VGND VGND VPWR VPWR OVHB\[6\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11626__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07929_ _07928_/Q _07952_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13544__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[13\].FF OVHB\[21\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[21\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ _10930_/CLK line[63] VGND VGND VPWR VPWR _10940_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08638__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10871_ _10870_/Q _10892_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12610_ _12638_/CLK line[58] VGND VGND VPWR VPWR _12610_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05062__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13590_ _13598_/CLK line[122] VGND VGND VPWR VPWR _13590_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ _12541_/A _12572_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05997__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[4\].TOBUF OVHB\[5\].VALID\[4\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08373__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[13\].VALID\[4\].FF OVHB\[13\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[13\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12472_ _12490_/CLK line[123] VGND VGND VPWR VPWR _12472_/Q sky130_fd_sc_hd__dfxtp_1
X_11423_ _11422_/Q _11452_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[8\].FF OVHB\[30\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[30\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07567__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11354_ _11370_/CLK line[124] VGND VGND VPWR VPWR _11354_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13719__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10305_ _10304_/Q _10332_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07286__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11285_ _11284_/Q _11312_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13024_ _13023_/Q _13027_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_10236_ _10248_/CLK line[125] VGND VGND VPWR VPWR _10236_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10143__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[13\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _06095_/CLK sky130_fd_sc_hd__clkbuf_4
X_10167_ _10166_/Q _10192_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05237__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10098_ _10100_/CLK line[62] VGND VGND VPWR VPWR _10098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13454__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08548__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13926_ A[5] VGND VGND VPWR VPWR _13934_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07452__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13857_ _13845_/CLK line[102] VGND VGND VPWR VPWR _13857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12808_ _12808_/A _12817_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13788_ _13787_/Q _13797_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12739_ _12741_/CLK line[103] VGND VGND VPWR VPWR _12739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11702__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09379__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06260_ _06244_/CLK line[85] VGND VGND VPWR VPWR _06260_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[9\].FF OVHB\[29\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[29\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08861__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05700__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05211_ _05210_/Q _05222_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10318__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].CGAND_A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06191_ _06190_/Q _06202_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__04940__A2_N _04940_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05142_ _05122_/CLK line[86] VGND VGND VPWR VPWR _05142_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].CGAND_A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13629__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12533__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05073_ _05072_/Q _05082_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_09950_ _09978_/CLK line[122] VGND VGND VPWR VPWR _09951_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[6\].FF OVHB\[11\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[11\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07627__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08901_ _08900_/Q _08932_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[20\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09881_ _09880_/Q _09912_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10053__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08832_ _08850_/CLK line[123] VGND VGND VPWR VPWR _08832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05975_ _05974_/Q _05992_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_08763_ _08763_/A _08792_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04926_ _04925_/X VGND VGND VPWR VPWR _04926_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07714_ _07724_/CLK line[124] VGND VGND VPWR VPWR _07714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04986__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08694_ _08710_/CLK line[60] VGND VGND VPWR VPWR _08694_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07362__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07645_ _07644_/Q _07672_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_07576_ _07572_/CLK line[61] VGND VGND VPWR VPWR _07576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06527_ _06526_/Q _06552_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_09315_ _09315_/CLK _09316_/X VGND VGND VPWR VPWR _09307_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12708__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09289__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08193__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06458_ _06464_/CLK line[62] VGND VGND VPWR VPWR _06458_/Q sky130_fd_sc_hd__dfxtp_1
X_09246_ _09352_/A wr VGND VGND VPWR VPWR _09246_/X sky130_fd_sc_hd__and2_1
XANTENNA__05610__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05409_ _05408_/Q _05432_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10228__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09177_ _09352_/A VGND VGND VPWR VPWR _09177_/Y sky130_fd_sc_hd__inv_2
X_06389_ _06388_/Q _06412_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08128_ _08134_/CLK line[48] VGND VGND VPWR VPWR _08128_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12443__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08059_ _08058_/Q _08092_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07537__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06441__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11070_ _11090_/CLK line[122] VGND VGND VPWR VPWR _11070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11059__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10021_ _10020_/Q _10052_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10541__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09752__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09107__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[9\].TOBUF OVHB\[3\].VALID\[9\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08368__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11972_ _11971_/Q _11977_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_13711_ _13701_/CLK line[35] VGND VGND VPWR VPWR _13711_/Q sky130_fd_sc_hd__dfxtp_1
X_10923_ _10903_/CLK line[41] VGND VGND VPWR VPWR _10924_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13642_ _13641_/Q _13657_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_10854_ _10853_/Q _10857_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12618__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _13559_/CLK line[100] VGND VGND VPWR VPWR _13573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ _10785_/CLK _10786_/X VGND VGND VPWR VPWR _10783_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _12523_/Q _12537_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06616__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12455_ _12449_/CLK line[101] VGND VGND VPWR VPWR _12455_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10716__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09927__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11406_ _11405_/Q _11417_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_12386_ _12385_/Q _12397_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_11337_ _11343_/CLK line[102] VGND VGND VPWR VPWR _11337_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06351__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11268_ _11267_/Q _11277_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13007_ _12999_/CLK line[97] VGND VGND VPWR VPWR _13007_/Q sky130_fd_sc_hd__dfxtp_1
X_10219_ _10217_/CLK line[103] VGND VGND VPWR VPWR _10220_/A sky130_fd_sc_hd__dfxtp_1
X_11199_ _11191_/CLK line[39] VGND VGND VPWR VPWR _11200_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13184__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13762__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08278__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05760_ _05756_/CLK line[127] VGND VGND VPWR VPWR _05761_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13481__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13909_ _13905_/X _13909_/B _13909_/C _13909_/D VGND VGND VPWR VPWR _13909_/X sky130_fd_sc_hd__and4b_4
X_05691_ _05690_/Q _05712_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_07430_ _07446_/CLK line[122] VGND VGND VPWR VPWR _07430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06376__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07361_ _07360_/Q _07392_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11432__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[4\].TOBUF OVHB\[10\].VALID\[4\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_09100_ _09099_/Q _09107_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_06312_ _06320_/CLK line[123] VGND VGND VPWR VPWR _06312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06526__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07292_ _07292_/CLK line[59] VGND VGND VPWR VPWR _07292_/Q sky130_fd_sc_hd__dfxtp_1
X_09031_ _09005_/CLK line[72] VGND VGND VPWR VPWR _09031_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10048__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06243_ _06243_/A _06272_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06174_ _06186_/CLK line[60] VGND VGND VPWR VPWR _06174_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08741__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13359__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05125_ _05125_/A _05152_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13937__A A[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09933_ _09925_/CLK line[100] VGND VGND VPWR VPWR _09933_/Q sky130_fd_sc_hd__dfxtp_1
X_05056_ _05058_/CLK line[61] VGND VGND VPWR VPWR _05056_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13656__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09864_ _09863_/Q _09877_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08815_ _08823_/CLK line[101] VGND VGND VPWR VPWR _08815_/Q sky130_fd_sc_hd__dfxtp_1
X_09795_ _09793_/CLK line[37] VGND VGND VPWR VPWR _09795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11607__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08746_ _08746_/A _08757_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07092__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05958_ _05984_/CLK line[80] VGND VGND VPWR VPWR _05958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08677_ _08663_/CLK line[38] VGND VGND VPWR VPWR _08677_/Q sky130_fd_sc_hd__dfxtp_1
X_05889_ _05889_/A _05922_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13822__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07628_ _07627_/Q _07637_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08916__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[0\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ _07539_/CLK line[39] VGND VGND VPWR VPWR _07559_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10570_ _10570_/A _10577_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09597__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05340__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09229_ _09241_/CLK line[34] VGND VGND VPWR VPWR _09229_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _12780_/CLK sky130_fd_sc_hd__clkbuf_4
X_12240_ _12240_/A _12257_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_12171_ _12177_/CLK line[99] VGND VGND VPWR VPWR _12171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12173__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07267__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[4\].VALID\[14\].TOBUF OVHB\[4\].VALID\[14\].FF/Q OVHB\[4\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_11122_ _11122_/A _11137_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11053_ _11063_/CLK line[100] VGND VGND VPWR VPWR _11053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09482__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10004_ _10003_/Q _10017_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10421__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05515__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DEC.DEC0.AND2_B A[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[1\].FF OVHB\[2\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[2\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11955_ _11945_/CLK line[15] VGND VGND VPWR VPWR _11955_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13732__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ _10905_/Q _10927_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11886_ _11885_/Q _11907_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07730__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12348__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13625_ _13631_/CLK line[10] VGND VGND VPWR VPWR _13625_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ _10843_/CLK line[1] VGND VGND VPWR VPWR _10837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[24\].VALID\[10\].TOBUF OVHB\[24\].VALID\[10\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_13556_ _13555_/Q _13587_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_10768_ _10767_/Q _10787_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
X_12507_ _12523_/CLK line[11] VGND VGND VPWR VPWR _12507_/Q sky130_fd_sc_hd__dfxtp_1
X_13487_ _13497_/CLK line[75] VGND VGND VPWR VPWR _13487_/Q sky130_fd_sc_hd__dfxtp_1
X_10699_ _10707_/CLK line[66] VGND VGND VPWR VPWR _10699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09657__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12438_ _12438_/A _12467_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12083__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12369_ _12387_/CLK line[76] VGND VGND VPWR VPWR _12369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06081__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[4\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _12395_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11277__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12811__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06930_ _06929_/Q _06937_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09392__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07905__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06861_ _06839_/CLK line[104] VGND VGND VPWR VPWR _06862_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08600_ _08600_/A _08617_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_05812_ _05811_/Q _05817_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_06792_ _06791_/Q _06797_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_09580_ _09580_/A _09597_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05743_ _05739_/CLK line[105] VGND VGND VPWR VPWR _05744_/A sky130_fd_sc_hd__dfxtp_1
X_08531_ _08541_/CLK line[99] VGND VGND VPWR VPWR _08532_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08462_ _08462_/A _08477_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_05674_ _05674_/A _05677_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07640__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07413_ _07393_/CLK line[100] VGND VGND VPWR VPWR _07413_/Q sky130_fd_sc_hd__dfxtp_1
X_08393_ _08383_/CLK line[36] VGND VGND VPWR VPWR _08393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12258__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11162__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07344_ _07343_/Q _07357_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06256__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[0\].VALID\[3\].FF OVHB\[0\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[0\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07275_ _07267_/CLK line[37] VGND VGND VPWR VPWR _07276_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09567__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06226_ _06225_/Q _06237_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_09014_ _09014_/A _09037_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08471__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13089__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06157_ _06147_/CLK line[38] VGND VGND VPWR VPWR _06158_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12571__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05108_ _05107_/Q _05117_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06088_ _06087_/Q _06097_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[13\].FF OVHB\[26\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[26\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12721__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09916_ _09915_/Q _09947_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_05039_ _05041_/CLK line[39] VGND VGND VPWR VPWR _05039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07815__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09847_ _09849_/CLK line[75] VGND VGND VPWR VPWR _09847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11337__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[3\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _12010_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_101_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09778_ _09778_/A _09807_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_08729_ _08749_/CLK line[76] VGND VGND VPWR VPWR _08729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[25\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11740_ _11739_/Q _11767_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08646__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11691_/CLK line[13] VGND VGND VPWR VPWR _11671_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11072__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13410_/CLK _13411_/X VGND VGND VPWR VPWR _13394_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ _10621_/Q _10647_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05070__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13272_/A wr VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__and2_1
X_10553_ _10571_/CLK line[14] VGND VGND VPWR VPWR _10553_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[4\].TOBUF OVHB\[17\].VALID\[4\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08381__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13272_ _13272_/A VGND VGND VPWR VPWR _13272_/Y sky130_fd_sc_hd__inv_2
X_10484_ _10483_/Q _10507_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12223_ _12227_/CLK line[0] VGND VGND VPWR VPWR _12223_/Q sky130_fd_sc_hd__dfxtp_1
X_12154_ _12153_/Q _12187_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[23\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _09350_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_97_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11105_ _11111_/CLK line[10] VGND VGND VPWR VPWR _11105_/Q sky130_fd_sc_hd__dfxtp_1
X_12085_ _12109_/CLK line[74] VGND VGND VPWR VPWR _12085_/Q sky130_fd_sc_hd__dfxtp_1
X_11036_ _11035_/Q _11067_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11247__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10151__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05245__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12987_ _12986_/Q _12992_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13462__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08556__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11938_ _11934_/CLK line[121] VGND VGND VPWR VPWR _11938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12078__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11869_ _11869_/A _11872_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_13608_ _13598_/CLK line[116] VGND VGND VPWR VPWR _13608_/Q sky130_fd_sc_hd__dfxtp_1
X_05390_ _05389_/Q _05397_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_13539_ _13539_/A _13552_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11710__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07060_ _07060_/A _07077_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06804__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06011_ _06023_/CLK line[99] VGND VGND VPWR VPWR _06011_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10326__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13637__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07962_ _07961_/Q _07987_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[23\].VALID\[3\].TOBUF OVHB\[23\].VALID\[3\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_09701_ _09632_/A wr VGND VGND VPWR VPWR _09701_/X sky130_fd_sc_hd__and2_1
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06913_ _06923_/CLK line[14] VGND VGND VPWR VPWR _06913_/Q sky130_fd_sc_hd__dfxtp_1
X_07893_ _07905_/CLK line[78] VGND VGND VPWR VPWR _07893_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _08965_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_56_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10061__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09632_ _09632_/A VGND VGND VPWR VPWR _09632_/Y sky130_fd_sc_hd__inv_2
X_06844_ _06844_/A _06867_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05155__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09563_ _09577_/CLK line[64] VGND VGND VPWR VPWR _09563_/Q sky130_fd_sc_hd__dfxtp_1
X_06775_ _06775_/CLK line[79] VGND VGND VPWR VPWR _06776_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08514_ _08513_/Q _08547_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04994__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05726_ _05725_/Q _05747_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09494_ _09493_/Q _09527_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07370__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _08473_/CLK line[74] VGND VGND VPWR VPWR _08445_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05657_ _05671_/CLK line[65] VGND VGND VPWR VPWR _05658_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _08375_/Q _08407_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
X_05588_ _05588_/A _05607_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[11\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07327_ _07327_/CLK line[75] VGND VGND VPWR VPWR _07328_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10086__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09297__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07258_ _07258_/A _07287_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[0\].FF OVHB\[25\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[25\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06209_ _06223_/CLK line[76] VGND VGND VPWR VPWR _06209_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10236__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07189_ _07183_/CLK line[12] VGND VGND VPWR VPWR _07190_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12451__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07545__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12910_ _12902_/CLK line[53] VGND VGND VPWR VPWR _12910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13890_ _13882_/CLK line[117] VGND VGND VPWR VPWR _13890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09760__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[15\].VALID\[9\].TOBUF OVHB\[15\].VALID\[9\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ _12840_/Q _12852_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ _12774_/CLK line[118] VGND VGND VPWR VPWR _12772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[30\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11723_ _11722_/Q _11732_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _05710_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11636_/CLK line[119] VGND VGND VPWR VPWR _11655_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[30\]_A1 _13459_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10605_ _10604_/Q _10612_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12626__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[22\].VALID\[11\].FF OVHB\[22\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[22\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11585_/A _11592_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13308_/CLK line[114] VGND VGND VPWR VPWR _13324_/Q sky130_fd_sc_hd__dfxtp_1
X_10536_ _10520_/CLK line[120] VGND VGND VPWR VPWR _10537_/A sky130_fd_sc_hd__dfxtp_1
X_13255_ _13255_/A _13272_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10467_ _10467_/A _10472_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09935__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12206_ _12204_/CLK line[115] VGND VGND VPWR VPWR _12207_/A sky130_fd_sc_hd__dfxtp_1
X_13186_ _13194_/CLK line[51] VGND VGND VPWR VPWR _13187_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10398_ _10384_/CLK line[57] VGND VGND VPWR VPWR _10398_/Q sky130_fd_sc_hd__dfxtp_1
X_12137_ _12136_/Q _12152_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[2\].FF OVHB\[23\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[23\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[24\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12068_ _12072_/CLK line[52] VGND VGND VPWR VPWR _12068_/Q sky130_fd_sc_hd__dfxtp_1
X_11019_ _11018_/Q _11032_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09670__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13192__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[12\].VALID\[13\].FF OVHB\[12\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[12\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08286__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06560_ _06560_/A _06587_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05511_ _05519_/CLK line[13] VGND VGND VPWR VPWR _05511_/Q sky130_fd_sc_hd__dfxtp_1
X_06491_ _06489_/CLK line[77] VGND VGND VPWR VPWR _06492_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05442_ _05441_/Q _05467_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_08230_ _08230_/CLK _08231_/X VGND VGND VPWR VPWR _08208_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_21_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[8\].TOBUF OVHB\[21\].VALID\[8\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_08161_ _13940_/X wr VGND VGND VPWR VPWR _08161_/X sky130_fd_sc_hd__and2_1
X_05373_ _05391_/CLK line[78] VGND VGND VPWR VPWR _05374_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[7\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11440__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07112_ _07111_/A VGND VGND VPWR VPWR _07112_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06534__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _05325_/CLK sky130_fd_sc_hd__clkbuf_4
X_08092_ _13940_/X VGND VGND VPWR VPWR _08092_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07043_ _07043_/CLK line[64] VGND VGND VPWR VPWR _07043_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[15\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09845__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06831__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13367__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08994_ _08972_/CLK line[55] VGND VGND VPWR VPWR _08995_/A sky130_fd_sc_hd__dfxtp_1
X_07945_ _07944_/Q _07952_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07876_ _07854_/CLK line[56] VGND VGND VPWR VPWR _07876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09615_ _09615_/A _09632_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06827_ _06827_/A _06832_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11615__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[29\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[4\].FF OVHB\[21\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[21\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06709__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09546_ _09554_/CLK line[51] VGND VGND VPWR VPWR _09546_/Q sky130_fd_sc_hd__dfxtp_1
X_06758_ _06740_/CLK line[57] VGND VGND VPWR VPWR _06758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05709_ _05709_/A _05712_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _09476_/Q _09492_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _06689_/A _06692_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ _08410_/CLK line[52] VGND VGND VPWR VPWR _08428_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08359_ _08358_/Q _08372_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[17\] _10873_/Z _07023_/Z _06533_/Z _05203_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[17] sky130_fd_sc_hd__mux4_1
XANTENNA_OVHB\[15\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11350__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].CG clk OVHB\[25\].CG/GATE VGND VGND VPWR VPWR OVHB\[25\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_11370_ _11370_/CLK line[117] VGND VGND VPWR VPWR _11371_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10321_ _10320_/Q _10332_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13040_ _13050_/CLK line[127] VGND VGND VPWR VPWR _13041_/A sky130_fd_sc_hd__dfxtp_1
X_10252_ _10248_/CLK line[118] VGND VGND VPWR VPWR _10252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13277__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12181__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10183_ _10183_/A _10192_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[14\].TOBUF OVHB\[17\].VALID\[14\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__07275__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[0\].TOBUF OVHB\[5\].VALID\[0\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13942_ _13944_/C _13946_/B _13944_/B _13944_/D VGND VGND VPWR VPWR _12151_/A sky130_fd_sc_hd__and4b_4
XFILLER_74_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13873_ _13872_/Q _13902_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11525__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12824_ _12820_/CLK line[28] VGND VGND VPWR VPWR _12824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[1\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05523__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12755_ _12754_/Q _12782_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13740__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[2\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/CLK line[29] VGND VGND VPWR VPWR _11706_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08834__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12686_ _12708_/CLK line[93] VGND VGND VPWR VPWR _12686_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12356__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11637_ _11637_/A _11662_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[10\].VALID\[13\].TOBUF OVHB\[10\].VALID\[13\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_128_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11568_ _11588_/CLK line[94] VGND VGND VPWR VPWR _11568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13307_ _13272_/A VGND VGND VPWR VPWR _13307_/Y sky130_fd_sc_hd__inv_2
X_10519_ _10519_/A _10542_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
X_11499_ _11498_/Q _11522_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
X_13238_ _13254_/CLK line[80] VGND VGND VPWR VPWR _13239_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12091__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10604__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13169_ _13169_/A _13202_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07185__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05991_ _13910_/X wr VGND VGND VPWR VPWR _05991_/X sky130_fd_sc_hd__and2_1
XFILLER_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _07724_/CLK line[117] VGND VGND VPWR VPWR _07730_/Q sky130_fd_sc_hd__dfxtp_1
X_04942_ _04921_/X _04931_/Y _04942_/C _04941_/X VGND VGND VPWR VPWR hit sky130_fd_sc_hd__and4_4
XANTENNA__07913__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07661_ _07660_/Q _07672_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09400_ _09414_/CLK line[127] VGND VGND VPWR VPWR _09400_/Q sky130_fd_sc_hd__dfxtp_1
X_06612_ _06596_/CLK line[118] VGND VGND VPWR VPWR _06612_/Q sky130_fd_sc_hd__dfxtp_1
X_07592_ _07572_/CLK line[54] VGND VGND VPWR VPWR _07592_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05433__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09331_ _09330_/Q _09352_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_06543_ _06542_/Q _06552_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09262_ _09256_/CLK line[49] VGND VGND VPWR VPWR _09262_/Q sky130_fd_sc_hd__dfxtp_1
X_06474_ _06464_/CLK line[55] VGND VGND VPWR VPWR _06475_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[7\].FF OVHB\[18\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[18\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08213_ _08212_/Q _08232_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12266__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05425_ _05424_/Q _05432_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_09193_ _09192_/Q _09212_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05356_ _05332_/CLK line[56] VGND VGND VPWR VPWR _05357_/A sky130_fd_sc_hd__dfxtp_1
X_08144_ _08134_/CLK line[50] VGND VGND VPWR VPWR _08144_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06264__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05287_ _05286_/Q _05292_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_08075_ _08074_/Q _08092_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[20\].INV _13965_/X VGND VGND VPWR VPWR OVHB\[20\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09575__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07026_ _07030_/CLK line[51] VGND VGND VPWR VPWR _07026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10514__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05608__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08977_ _08977_/A _09002_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[20\]_A0 _10039_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07928_ _07946_/CLK line[94] VGND VGND VPWR VPWR _07928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07823__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07859_ _07858_/Q _07882_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06439__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10870_ _10872_/CLK line[31] VGND VGND VPWR VPWR _10870_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[13\].TOBUF OVHB\[30\].VALID\[13\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05921__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ _09528_/Q _09562_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ _12560_/CLK line[26] VGND VGND VPWR VPWR _12541_/A sky130_fd_sc_hd__dfxtp_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12470_/Q _12502_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11080__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[3\].VALID\[5\].TOBUF OVHB\[3\].VALID\[5\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06174__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11422_ _11440_/CLK line[27] VGND VGND VPWR VPWR _11422_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[8\].TOBUF OVHB\[28\].VALID\[8\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12904__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11353_ _11352_/Q _11382_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10304_ _10314_/CLK line[28] VGND VGND VPWR VPWR _10304_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[9\].FF OVHB\[16\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[16\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11284_ _11302_/CLK line[92] VGND VGND VPWR VPWR _11284_/Q sky130_fd_sc_hd__dfxtp_1
X_13023_ _12999_/CLK line[105] VGND VGND VPWR VPWR _13023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[20\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10235_ _10235_/A _10262_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10166_ _10188_/CLK line[93] VGND VGND VPWR VPWR _10166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10097_ _10096_/Q _10122_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13925_ A[4] VGND VGND VPWR VPWR _13933_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_OVHB\[13\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11255__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13856_ _13856_/A _13867_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06349__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05253__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12807_ _12803_/CLK line[6] VGND VGND VPWR VPWR _12808_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13787_ _13763_/CLK line[70] VGND VGND VPWR VPWR _13787_/Q sky130_fd_sc_hd__dfxtp_1
X_10999_ _10998_/Q _11032_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13470__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12738_ _12737_/Q _12747_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08564__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _12667_/CLK line[71] VGND VGND VPWR VPWR _12669_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08861__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05210_ _05214_/CLK line[117] VGND VGND VPWR VPWR _05210_/Q sky130_fd_sc_hd__dfxtp_1
X_06190_ _06186_/CLK line[53] VGND VGND VPWR VPWR _06190_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05141_ _05140_/Q _05152_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].V OVHB\[3\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[3\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_DATA\[0\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05072_ _05058_/CLK line[54] VGND VGND VPWR VPWR _05072_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06812__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].CGAND_A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08900_ _08922_/CLK line[26] VGND VGND VPWR VPWR _08900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09880_ _09908_/CLK line[90] VGND VGND VPWR VPWR _09880_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05428__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[0\].TOBUF OVHB\[10\].VALID\[0\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_08831_ _08830_/Q _08862_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13645__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08739__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08762_ _08762_/CLK line[91] VGND VGND VPWR VPWR _08763_/A sky130_fd_sc_hd__dfxtp_1
X_05974_ _05984_/CLK line[82] VGND VGND VPWR VPWR _05974_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[13\].FF OVHB\[3\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[3\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07713_ _07712_/Q _07742_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
X_04925_ A_h[15] _04924_/Y _04922_/Y _04923_/B VGND VGND VPWR VPWR _04925_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08693_ _08693_/A _08722_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07644_ _07644_/CLK line[92] VGND VGND VPWR VPWR _07644_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05163__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07575_ _07574_/Q _07602_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13380__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09314_ _09313_/Q _09317_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_06526_ _06528_/CLK line[93] VGND VGND VPWR VPWR _06526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09245_ _09245_/CLK _09246_/X VGND VGND VPWR VPWR _09241_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_90_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06457_ _06457_/A _06482_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _08265_/CLK sky130_fd_sc_hd__clkbuf_4
X_05408_ _05424_/CLK line[94] VGND VGND VPWR VPWR _05408_/Q sky130_fd_sc_hd__dfxtp_1
X_09176_ _09352_/A wr VGND VGND VPWR VPWR _09176_/X sky130_fd_sc_hd__and2_1
X_06388_ _06408_/CLK line[30] VGND VGND VPWR VPWR _06388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08127_ _13940_/X VGND VGND VPWR VPWR _08127_/Y sky130_fd_sc_hd__inv_2
X_05339_ _05338_/Q _05362_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08058_ _08070_/CLK line[16] VGND VGND VPWR VPWR _08058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07009_ _07008_/Q _07042_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10244__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[31\].VOBUF OVHB\[31\].V/Q OVHB\[31\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__10822__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05338__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10020_ _10042_/CLK line[26] VGND VGND VPWR VPWR _10020_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10541__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13555__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07553__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[31\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _11835_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_17_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11971_ _11945_/CLK line[8] VGND VGND VPWR VPWR _11971_/Q sky130_fd_sc_hd__dfxtp_1
X_13710_ _13709_/Q _13727_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10922_ _10921_/Q _10927_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[11\].FF OVHB\[27\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[27\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13641_ _13631_/CLK line[3] VGND VGND VPWR VPWR _13641_/Q sky130_fd_sc_hd__dfxtp_1
X_10853_ _10843_/CLK line[9] VGND VGND VPWR VPWR _10853_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[10\].TOBUF OVHB\[4\].VALID\[10\].FF/Q OVHB\[4\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11803__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _13571_/Q _13587_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_10784_ _10783_/Q _10787_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05801__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _12523_/CLK line[4] VGND VGND VPWR VPWR _12523_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10419__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12454_ _12453_/Q _12467_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06482__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10716__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11405_ _11395_/CLK line[5] VGND VGND VPWR VPWR _11405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12634__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _12387_/CLK line[69] VGND VGND VPWR VPWR _12385_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[0\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _05080_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07728__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11336_ _11336_/A _11347_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[2\].FF OVHB\[9\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[9\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11267_ _11251_/CLK line[70] VGND VGND VPWR VPWR _11267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09943__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13006_ _13005_/Q _13027_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_10218_ _10218_/A _10227_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11198_ _11197_/Q _11207_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[21\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[13\].FF OVHB\[17\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[17\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10149_ _10145_/CLK line[71] VGND VGND VPWR VPWR _10149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07463__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06079__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _13905_/X _13909_/C _13909_/B _13909_/D VGND VGND VPWR VPWR _13908_/X sky130_fd_sc_hd__and4bb_4
X_05690_ _05708_/CLK line[95] VGND VGND VPWR VPWR _05690_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06657__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12809__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13839_ _13845_/CLK line[108] VGND VGND VPWR VPWR _13839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[2\]_A0 _09160_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06376__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _11450_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08294__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07360_ _07380_/CLK line[90] VGND VGND VPWR VPWR _07360_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06311_ _06311_/A _06342_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[20\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _08580_/CLK sky130_fd_sc_hd__clkbuf_4
X_07291_ _07290_/Q _07322_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_09030_ _09030_/A _09037_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_06242_ _06244_/CLK line[91] VGND VGND VPWR VPWR _06243_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].INV _13988_/X VGND VGND VPWR VPWR OVHB\[5\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12544__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06173_ _06172_/Q _06202_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07638__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05124_ _05122_/CLK line[92] VGND VGND VPWR VPWR _05125_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06542__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09932_ _09932_/A _09947_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_05055_ _05054_/Q _05082_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09853__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09863_ _09849_/CLK line[68] VGND VGND VPWR VPWR _09863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08814_ _08813_/Q _08827_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08469__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09794_ _09793_/Q _09807_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07951__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08745_ _08749_/CLK line[69] VGND VGND VPWR VPWR _08746_/A sky130_fd_sc_hd__dfxtp_1
X_05957_ _13910_/X VGND VGND VPWR VPWR _05957_/Y sky130_fd_sc_hd__inv_2
XOVHB\[7\].VALID\[4\].FF OVHB\[7\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[7\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08676_ _08675_/Q _08687_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_05888_ _05902_/CLK line[48] VGND VGND VPWR VPWR _05889_/A sky130_fd_sc_hd__dfxtp_1
X_07627_ _07633_/CLK line[70] VGND VGND VPWR VPWR _07627_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12719__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07558_ _07557_/Q _07567_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06509_ _06489_/CLK line[71] VGND VGND VPWR VPWR _06509_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[12\].TOBUF OVHB\[27\].VALID\[12\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_07489_ _07467_/CLK line[7] VGND VGND VPWR VPWR _07489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09228_ _09228_/A _09247_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09159_ _09147_/CLK line[2] VGND VGND VPWR VPWR _09159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06452__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _12169_/Q _12187_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11121_ _11111_/CLK line[3] VGND VGND VPWR VPWR _11122_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05068__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11052_ _11051_/Q _11067_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08022__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13285__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10003_ _10011_/CLK line[4] VGND VGND VPWR VPWR _10003_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08379__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07283__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[17\].VALID\[0\].TOBUF OVHB\[17\].VALID\[0\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ _11953_/Q _11977_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[11\].TOBUF OVHB\[20\].VALID\[11\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10905_ _10903_/CLK line[47] VGND VGND VPWR VPWR _10905_/Q sky130_fd_sc_hd__dfxtp_1
X_11885_ _11901_/CLK line[111] VGND VGND VPWR VPWR _11885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11533__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13624_ _13624_/A _13657_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06627__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10836_ _10835_/Q _10857_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05531__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09003__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[6\].FF OVHB\[5\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[5\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13555_ _13559_/CLK line[106] VGND VGND VPWR VPWR _13555_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10149__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10767_ _10783_/CLK line[97] VGND VGND VPWR VPWR _10767_/Q sky130_fd_sc_hd__dfxtp_1
X_12506_ _12505_/Q _12537_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08842__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _13485_/Q _13517_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_10698_ _10697_/Q _10717_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_12437_ _12449_/CLK line[107] VGND VGND VPWR VPWR _12438_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07458__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12368_ _12368_/A _12397_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11319_ _11343_/CLK line[108] VGND VGND VPWR VPWR _11319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12299_ _12311_/CLK line[44] VGND VGND VPWR VPWR _12299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11708__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06860_ _06860_/A _06867_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07193__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05706__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05811_ _05799_/CLK line[8] VGND VGND VPWR VPWR _05811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06791_ _06775_/CLK line[72] VGND VGND VPWR VPWR _06791_/Q sky130_fd_sc_hd__dfxtp_1
X_08530_ _08530_/A _08547_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05742_ _05741_/Q _05747_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05291__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08461_ _08473_/CLK line[67] VGND VGND VPWR VPWR _08462_/A sky130_fd_sc_hd__dfxtp_1
X_05673_ _05671_/CLK line[73] VGND VGND VPWR VPWR _05674_/A sky130_fd_sc_hd__dfxtp_1
X_07412_ _07411_/Q _07427_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08392_ _08391_/Q _08407_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05441__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10059__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07343_ _07327_/CLK line[68] VGND VGND VPWR VPWR _07343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07274_ _07273_/Q _07287_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[20\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09013_ _09005_/CLK line[78] VGND VGND VPWR VPWR _09014_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13948__A A_h[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06225_ _06223_/CLK line[69] VGND VGND VPWR VPWR _06225_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12274__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12852__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[11\].FF OVHB\[13\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[13\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07368__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06156_ _06155_/Q _06167_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[8\].FF OVHB\[3\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[3\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12571__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05107_ _05093_/CLK line[70] VGND VGND VPWR VPWR _05107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06087_ _06077_/CLK line[6] VGND VGND VPWR VPWR _06087_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09583__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05466__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09915_ _09925_/CLK line[106] VGND VGND VPWR VPWR _09915_/Q sky130_fd_sc_hd__dfxtp_1
X_05038_ _05037_/Q _05047_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10522__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09846_ _09845_/Q _09877_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05616__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09777_ _09793_/CLK line[43] VGND VGND VPWR VPWR _09778_/A sky130_fd_sc_hd__dfxtp_1
X_06989_ _07001_/CLK line[34] VGND VGND VPWR VPWR _06990_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13833__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08728_ _08727_/Q _08757_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07831__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12449__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08659_ _08663_/CLK line[44] VGND VGND VPWR VPWR _08659_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11669_/Q _11697_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10627_/CLK line[45] VGND VGND VPWR VPWR _10621_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13340_/CLK _13341_/X VGND VGND VPWR VPWR _13308_/CLK sky130_fd_sc_hd__dlclkp_1
X_10552_ _10551_/Q _10577_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13271_ _13272_/A wr VGND VGND VPWR VPWR _13271_/X sky130_fd_sc_hd__and2_1
XOVHB\[15\].VALID\[5\].TOBUF OVHB\[15\].VALID\[5\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_10483_ _10473_/CLK line[110] VGND VGND VPWR VPWR _10483_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[2\].FF OVHB\[31\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[31\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06182__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12222_ _12151_/A VGND VGND VPWR VPWR _12222_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12153_ _12177_/CLK line[96] VGND VGND VPWR VPWR _12153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12912__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09493__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11104_ _11103_/Q _11137_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12084_ _12084_/A _12117_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11035_ _11063_/CLK line[106] VGND VGND VPWR VPWR _11035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08687__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[9\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12986_ _12962_/CLK line[88] VGND VGND VPWR VPWR _12986_/Q sky130_fd_sc_hd__dfxtp_1
X_11937_ _11936_/Q _11942_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[3\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11263__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06357__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11868_ _11846_/CLK line[89] VGND VGND VPWR VPWR _11869_/A sky130_fd_sc_hd__dfxtp_1
X_10819_ _10818_/Q _10822_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_13607_ _13606_/Q _13622_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_11799_ _11799_/A _11802_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09668__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08572__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13538_ _13528_/CLK line[84] VGND VGND VPWR VPWR _13539_/A sky130_fd_sc_hd__dfxtp_1
X_13469_ _13468_/Q _13482_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06010_ _06009_/Q _06027_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12822__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[13\].FF OVHB\[8\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[8\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10192__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[12\].VALID\[0\].FF OVHB\[12\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[12\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06820__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09981__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07961_ _07981_/CLK line[109] VGND VGND VPWR VPWR _07961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11438__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09700_ _09700_/CLK _09701_/X VGND VGND VPWR VPWR _09694_/CLK sky130_fd_sc_hd__dlclkp_1
X_06912_ _06911_/Q _06937_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07892_ _07891_/Q _07917_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[4\].TOBUF OVHB\[21\].VALID\[4\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_09631_ _09632_/A wr VGND VGND VPWR VPWR _09631_/X sky130_fd_sc_hd__and2_1
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06843_ _06839_/CLK line[110] VGND VGND VPWR VPWR _06844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13653__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09562_ _09632_/A VGND VGND VPWR VPWR _09562_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08747__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06774_ _06773_/Q _06797_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_08513_ _08541_/CLK line[96] VGND VGND VPWR VPWR _08513_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07006__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05725_ _05739_/CLK line[111] VGND VGND VPWR VPWR _05725_/Q sky130_fd_sc_hd__dfxtp_1
X_09493_ _09507_/CLK line[32] VGND VGND VPWR VPWR _09493_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11173__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _08443_/Q _08477_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_05656_ _05655_/Q _05677_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05171__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _08383_/CLK line[42] VGND VGND VPWR VPWR _08375_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10367__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05587_ _05575_/CLK line[33] VGND VGND VPWR VPWR _05588_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11901__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07326_ _07325_/Q _07357_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08482__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10086__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07257_ _07267_/CLK line[43] VGND VGND VPWR VPWR _07258_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07098__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06208_ _06207_/Q _06237_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07188_ _07187_/Q _07217_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13828__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06139_ _06147_/CLK line[44] VGND VGND VPWR VPWR _06140_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[5\].FF OVHB\[28\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[28\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06730__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11348__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10252__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05346__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09829_ _09829_/A _09842_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13563__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12840_ _12820_/CLK line[21] VGND VGND VPWR VPWR _12840_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[2\].FF OVHB\[10\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[10\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08657__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07561__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12179__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _12770_/Q _12782_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11661__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11722_ _11706_/CLK line[22] VGND VGND VPWR VPWR _11722_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[10\].TOBUF OVHB\[17\].VALID\[10\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_11653_ _11653_/A _11662_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_MUX.MUX\[30\]_A2 _09609_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11811__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09488__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTIE VGND VGND VPWR VPWR TIE/HI TIE/LO sky130_fd_sc_hd__conb_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _10594_/CLK line[23] VGND VGND VPWR VPWR _10604_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06905__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ _11588_/CLK line[87] VGND VGND VPWR VPWR _11585_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13323_ _13322_/Q _13342_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10427__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ _10535_/A _10542_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13254_ _13254_/CLK line[82] VGND VGND VPWR VPWR _13255_/A sky130_fd_sc_hd__dfxtp_1
X_10466_ _10466_/CLK line[88] VGND VGND VPWR VPWR _10467_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13738__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ _12204_/Q _12222_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_13185_ _13184_/Q _13202_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_10397_ _10396_/Q _10402_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07736__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _12130_/CLK line[83] VGND VGND VPWR VPWR _12136_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04939__A1_N A_h[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11836__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10162__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ _12066_/Q _12082_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11018_ _11002_/CLK line[84] VGND VGND VPWR VPWR _11018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07471__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[7\].FF OVHB\[26\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[26\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12089__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12969_ _12969_/A _12992_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_05510_ _05509_/Q _05537_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06087__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06490_ _06489_/Q _06517_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05441_ _05445_/CLK line[109] VGND VGND VPWR VPWR _05441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09398__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08160_ _08160_/CLK _08161_/X VGND VGND VPWR VPWR _08134_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_119_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05372_ _05371_/Q _05397_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
X_07111_ _07111_/A wr VGND VGND VPWR VPWR _07111_/X sky130_fd_sc_hd__and2_1
XANTENNA__10337__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08091_ _13940_/X wr VGND VGND VPWR VPWR _08091_/X sky130_fd_sc_hd__and2_1
XANTENNA__07496__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07042_ _07111_/A VGND VGND VPWR VPWR _07042_/Y sky130_fd_sc_hd__inv_2
XANTENNA_MUX.MUX\[15\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12552__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07646__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08993_ _08993_/A _09002_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11168__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07944_ _07946_/CLK line[87] VGND VGND VPWR VPWR _07944_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[9\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09861__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07875_ _07875_/A _07882_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_09614_ _09626_/CLK line[82] VGND VGND VPWR VPWR _09615_/A sky130_fd_sc_hd__dfxtp_1
X_06826_ _06802_/CLK line[88] VGND VGND VPWR VPWR _06827_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10800__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09545_ _09544_/Q _09562_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06757_ _06756_/Q _06762_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05708_ _05708_/CLK line[89] VGND VGND VPWR VPWR _05709_/A sky130_fd_sc_hd__dfxtp_1
X_09476_ _09482_/CLK line[19] VGND VGND VPWR VPWR _09476_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ _06682_/CLK line[25] VGND VGND VPWR VPWR _06689_/A sky130_fd_sc_hd__dfxtp_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _08426_/Q _08442_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12727__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05639_ _05639_/A _05642_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[9\].FF OVHB\[24\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[24\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _08358_/CLK line[20] VGND VGND VPWR VPWR _08358_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[11\].FF OVHB\[4\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[4\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09101__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07309_ _07309_/A _07322_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_08289_ _08288_/Q _08302_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13201__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10320_ _10314_/CLK line[21] VGND VGND VPWR VPWR _10320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10251_ _10250_/Q _10262_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06460__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10182_ _10188_/CLK line[86] VGND VGND VPWR VPWR _10183_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11078__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05076__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13941_ _13944_/C _13944_/B _13946_/B _13944_/D VGND VGND VPWR VPWR _11311_/A sky130_fd_sc_hd__and4bb_4
XOVHB\[3\].VALID\[1\].TOBUF OVHB\[3\].VALID\[1\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13293__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08387__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13872_ _13882_/CLK line[123] VGND VGND VPWR VPWR _13872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[4\].TOBUF OVHB\[28\].VALID\[4\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12823_ _12822_/Q _12852_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12774_/CLK line[124] VGND VGND VPWR VPWR _12754_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11705_ _11704_/Q _11732_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VOBUF OVHB\[26\].V/Q OVHB\[26\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12684_/Q _12712_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06635__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11636_ _11636_/CLK line[125] VGND VGND VPWR VPWR _11637_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09011__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _11566_/Q _11592_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_13306_ _13272_/A wr VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__and2_1
XANTENNA__08850__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10518_ _10520_/CLK line[126] VGND VGND VPWR VPWR _10519_/A sky130_fd_sc_hd__dfxtp_1
X_11498_ _11500_/CLK line[62] VGND VGND VPWR VPWR _11498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13468__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13237_ _13272_/A VGND VGND VPWR VPWR _13237_/Y sky130_fd_sc_hd__inv_2
X_10449_ _10448_/Q _10472_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13168_ _13194_/CLK line[48] VGND VGND VPWR VPWR _13169_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12119_ _12118_/Q _12152_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13099_ _13098_/Q _13132_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_05990_ _05990_/CLK _05991_/X VGND VGND VPWR VPWR _05984_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09036__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04941_ _04937_/X _04938_/X _04941_/C _04940_/X VGND VGND VPWR VPWR _04941_/X sky130_fd_sc_hd__and4_4
XFILLER_133_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11716__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07660_ _07644_/CLK line[85] VGND VGND VPWR VPWR _07660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06611_ _06611_/A _06622_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[21\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07591_ _07590_/Q _07602_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12397__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09330_ _09320_/CLK line[95] VGND VGND VPWR VPWR _09330_/Q sky130_fd_sc_hd__dfxtp_1
X_06542_ _06528_/CLK line[86] VGND VGND VPWR VPWR _06542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09261_ _09260_/Q _09282_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[11\].FF OVHB\[18\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[18\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06473_ _06472_/Q _06482_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_08212_ _08208_/CLK line[81] VGND VGND VPWR VPWR _08212_/Q sky130_fd_sc_hd__dfxtp_1
X_05424_ _05424_/CLK line[87] VGND VGND VPWR VPWR _05424_/Q sky130_fd_sc_hd__dfxtp_1
X_09192_ _09200_/CLK line[17] VGND VGND VPWR VPWR _09192_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10067__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08143_ _08143_/A _08162_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_05355_ _05354_/Q _05362_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08760__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08074_ _08070_/CLK line[18] VGND VGND VPWR VPWR _08074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05286_ _05278_/CLK line[24] VGND VGND VPWR VPWR _05286_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13378__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07025_ _07024_/Q _07042_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12282__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07376__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08976_ _08972_/CLK line[61] VGND VGND VPWR VPWR _08977_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09591__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[20\]_A1 _13469_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07927_ _07926_/Q _07952_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[11\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13691__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10530__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07858_ _07854_/CLK line[62] VGND VGND VPWR VPWR _07858_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05624__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06809_ _06808_/Q _06832_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08000__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07789_ _07788_/Q _07812_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13841__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08935__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05921__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09528_ _09554_/CLK line[48] VGND VGND VPWR VPWR _09528_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09459_ _09458_/Q _09492_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12470_ _12490_/CLK line[122] VGND VGND VPWR VPWR _12470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[30\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11421_ _11420_/Q _11452_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09766__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[6\].TOBUF OVHB\[1\].VALID\[6\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_11352_ _11370_/CLK line[123] VGND VGND VPWR VPWR _11352_/Q sky130_fd_sc_hd__dfxtp_1
X_10303_ _10302_/Q _10332_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13866__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10705__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12192__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[9\].TOBUF OVHB\[26\].VALID\[9\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_11283_ _11283_/A _11312_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06190__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ _13021_/Q _13027_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_10234_ _10248_/CLK line[124] VGND VGND VPWR VPWR _10235_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10165_ _10164_/Q _10192_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10096_ _10100_/CLK line[61] VGND VGND VPWR VPWR _10096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10440__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _13922_/B _13923_/B _13923_/C _13923_/D VGND VGND VPWR VPWR _09352_/A sky130_fd_sc_hd__and4_4
XFILLER_63_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _13845_/CLK line[101] VGND VGND VPWR VPWR _13856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ _12805_/Q _12817_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_10998_ _11002_/CLK line[80] VGND VGND VPWR VPWR _10998_/Q sky130_fd_sc_hd__dfxtp_1
X_13786_ _13785_/Q _13797_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12367__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[27\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12737_ _12741_/CLK line[102] VGND VGND VPWR VPWR _12737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11271__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06365__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _12667_/Q _12677_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11619_ _11605_/CLK line[103] VGND VGND VPWR VPWR _11619_/Q sky130_fd_sc_hd__dfxtp_1
X_12599_ _12601_/CLK line[39] VGND VGND VPWR VPWR _12599_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09676__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05140_ _05122_/CLK line[85] VGND VGND VPWR VPWR _05140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13198__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10615__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05071_ _05070_/Q _05082_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08830_ _08850_/CLK line[122] VGND VGND VPWR VPWR _08830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12830__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].CGAND_A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07924__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08761_ _08760_/Q _08792_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05973_ _05972_/Q _05992_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11446__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07712_ _07724_/CLK line[123] VGND VGND VPWR VPWR _07712_/Q sky130_fd_sc_hd__dfxtp_1
X_04924_ _04924_/A VGND VGND VPWR VPWR _04924_/Y sky130_fd_sc_hd__inv_2
XOVHB\[15\].CG clk OVHB\[15\].CGAND/X VGND VGND VPWR VPWR OVHB\[15\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_08692_ _08710_/CLK line[59] VGND VGND VPWR VPWR _08693_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07643_ _07642_/Q _07672_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_07574_ _07572_/CLK line[60] VGND VGND VPWR VPWR _07574_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[12\].TOBUF OVHB\[7\].VALID\[12\].FF/Q OVHB\[7\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09313_ _09307_/CLK line[73] VGND VGND VPWR VPWR _09313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06525_ _06524_/Q _06552_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11181__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09244_ _09244_/A _09247_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06275__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06456_ _06464_/CLK line[61] VGND VGND VPWR VPWR _06457_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05407_ _05406_/Q _05432_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_09175_ _09175_/CLK _09176_/X VGND VGND VPWR VPWR _09147_/CLK sky130_fd_sc_hd__dlclkp_1
X_06387_ _06386_/Q _06412_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08126_ _13940_/X wr VGND VGND VPWR VPWR _08126_/X sky130_fd_sc_hd__and2_1
XANTENNA__08490__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05338_ _05332_/CLK line[62] VGND VGND VPWR VPWR _05338_/Q sky130_fd_sc_hd__dfxtp_1
X_08057_ _13940_/X VGND VGND VPWR VPWR _08057_/Y sky130_fd_sc_hd__inv_2
X_05269_ _05268_/Q _05292_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[0\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07008_ _07030_/CLK line[48] VGND VGND VPWR VPWR _07008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[0\].VALID\[11\].TOBUF OVHB\[0\].VALID\[11\].FF/Q OVHB\[0\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_08959_ _08947_/CLK line[39] VGND VGND VPWR VPWR _08960_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DEC.DEC0.AND2_A_N A[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11356__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[28\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11970_ _11970_/A _11977_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05354__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10921_ _10903_/CLK line[40] VGND VGND VPWR VPWR _10921_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13571__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08665__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13640_ _13639_/Q _13657_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10852_ _10851_/Q _10857_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ _10783_/CLK line[105] VGND VGND VPWR VPWR _10783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _13559_/CLK line[99] VGND VGND VPWR VPWR _13571_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12521_/Q _12537_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12453_ _12449_/CLK line[100] VGND VGND VPWR VPWR _12453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06913__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11404_ _11404_/A _11417_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_12384_ _12383_/Q _12397_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11335_ _11343_/CLK line[101] VGND VGND VPWR VPWR _11336_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[1\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05529__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11266_ _11265_/Q _11277_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13746__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10217_ _10217_/CLK line[102] VGND VGND VPWR VPWR _10218_/A sky130_fd_sc_hd__dfxtp_1
X_13005_ _12999_/CLK line[111] VGND VGND VPWR VPWR _13005_/Q sky130_fd_sc_hd__dfxtp_1
X_11197_ _11191_/CLK line[38] VGND VGND VPWR VPWR _11197_/Q sky130_fd_sc_hd__dfxtp_1
X_10148_ _10148_/A _10157_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10170__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10079_ _10073_/CLK line[39] VGND VGND VPWR VPWR _10080_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05264__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13907_ _13905_/X _13909_/B _13909_/C _13909_/D VGND VGND VPWR VPWR _13907_/X sky130_fd_sc_hd__and4bb_4
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[18\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13838_ _13837_/Q _13867_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[2\]_A1 _05030_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12097__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13769_ _13763_/CLK line[76] VGND VGND VPWR VPWR _13769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06310_ _06320_/CLK line[122] VGND VGND VPWR VPWR _06311_/A sky130_fd_sc_hd__dfxtp_1
X_07290_ _07292_/CLK line[58] VGND VGND VPWR VPWR _07290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_MUX.MUX\[10\]_A0 _11386_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06241_ _06240_/Q _06272_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06172_ _06186_/CLK line[59] VGND VGND VPWR VPWR _06172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[19\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _07950_/CLK sky130_fd_sc_hd__clkbuf_4
X_05123_ _05122_/Q _05152_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10345__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[8\].VALID\[6\].TOBUF OVHB\[8\].VALID\[6\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__05439__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09931_ _09925_/CLK line[99] VGND VGND VPWR VPWR _09932_/A sky130_fd_sc_hd__dfxtp_1
X_05054_ _05058_/CLK line[60] VGND VGND VPWR VPWR _05054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12560__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09862_ _09861_/Q _09877_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07654__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08813_ _08823_/CLK line[100] VGND VGND VPWR VPWR _08813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09793_ _09793_/CLK line[36] VGND VGND VPWR VPWR _09793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05956_ _13910_/X wr VGND VGND VPWR VPWR _05956_/X sky130_fd_sc_hd__and2_1
X_08744_ _08743_/Q _08757_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07951__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08675_ _08663_/CLK line[37] VGND VGND VPWR VPWR _08675_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[13\].TOBUF OVHB\[23\].VALID\[13\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_22_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05887_ _13910_/X VGND VGND VPWR VPWR _05887_/Y sky130_fd_sc_hd__inv_2
XOVHB\[9\].VALID\[11\].FF OVHB\[9\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[9\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07626_ _07625_/Q _07637_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05902__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ _07539_/CLK line[38] VGND VGND VPWR VPWR _07557_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06508_ _06507_/Q _06517_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
X_07488_ _07487_/Q _07497_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_09227_ _09241_/CLK line[33] VGND VGND VPWR VPWR _09228_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12735__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06439_ _06421_/CLK line[39] VGND VGND VPWR VPWR _06440_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07829__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09158_ _09157_/Q _09177_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_08109_ _08113_/CLK line[34] VGND VGND VPWR VPWR _08109_/Q sky130_fd_sc_hd__dfxtp_1
X_09089_ _09085_/CLK line[98] VGND VGND VPWR VPWR _09089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11120_ _11119_/Q _11137_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11051_ _11063_/CLK line[99] VGND VGND VPWR VPWR _11051_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12470__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[18\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _07565_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[30\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10002_ _10001_/Q _10017_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11086__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[15\].VALID\[1\].TOBUF OVHB\[15\].VALID\[1\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11953_ _11945_/CLK line[14] VGND VGND VPWR VPWR _11953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08395__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10904_ _10903_/Q _10927_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11884_ _11883_/Q _11907_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_13623_ _13631_/CLK line[0] VGND VGND VPWR VPWR _13624_/A sky130_fd_sc_hd__dfxtp_1
X_10835_ _10843_/CLK line[15] VGND VGND VPWR VPWR _10835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13554_ _13553_/Q _13587_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_10766_ _10765_/Q _10787_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12505_ _12523_/CLK line[10] VGND VGND VPWR VPWR _12505_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12645__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10697_ _10707_/CLK line[65] VGND VGND VPWR VPWR _10697_/Q sky130_fd_sc_hd__dfxtp_1
X_13485_ _13497_/CLK line[74] VGND VGND VPWR VPWR _13485_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[0\].FF OVHB\[20\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[20\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06643__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12436_ _12435_/Q _12467_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_12367_ _12387_/CLK line[75] VGND VGND VPWR VPWR _12368_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09954__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11318_ _11317_/Q _11347_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_12298_ _12298_/A _12327_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13476__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11249_ _11251_/CLK line[76] VGND VGND VPWR VPWR _11250_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05810_ _05810_/A _05817_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_06790_ _06789_/Q _06797_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05572__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05741_ _05739_/CLK line[104] VGND VGND VPWR VPWR _05741_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11724__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ _08459_/Q _08477_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05291__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05672_ _05671_/Q _05677_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06818__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07411_ _07393_/CLK line[99] VGND VGND VPWR VPWR _07411_/Q sky130_fd_sc_hd__dfxtp_1
X_08391_ _08383_/CLK line[35] VGND VGND VPWR VPWR _08391_/Q sky130_fd_sc_hd__dfxtp_1
X_07342_ _07341_/Q _07357_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[19\].VALID\[1\].FF OVHB\[19\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[19\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[0\].TOBUF OVHB\[21\].VALID\[0\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_07273_ _07267_/CLK line[36] VGND VGND VPWR VPWR _07273_/Q sky130_fd_sc_hd__dfxtp_1
X_09012_ _09011_/Q _09037_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
X_06224_ _06223_/Q _06237_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06553__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10075__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06155_ _06147_/CLK line[37] VGND VGND VPWR VPWR _06155_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05169__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05106_ _05105_/Q _05117_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05747__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06086_ _06086_/A _06097_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13386__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09914_ _09913_/Q _09947_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05466__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05037_ _05041_/CLK line[38] VGND VGND VPWR VPWR _05037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07384__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09845_ _09849_/CLK line[74] VGND VGND VPWR VPWR _09845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09776_ _09775_/Q _09807_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
X_06988_ _06987_/Q _07007_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_08727_ _08749_/CLK line[75] VGND VGND VPWR VPWR _08727_/Q sky130_fd_sc_hd__dfxtp_1
X_05939_ _05929_/CLK line[66] VGND VGND VPWR VPWR _05939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11634__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06728__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08658_ _08657_/Q _08687_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05632__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07633_/CLK line[76] VGND VGND VPWR VPWR _07610_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08609_/CLK line[12] VGND VGND VPWR VPWR _08589_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08943__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10620_ _10619_/Q _10647_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _10571_/CLK line[13] VGND VGND VPWR VPWR _10551_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07559__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10482_ _10481_/Q _10507_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_13270_ _13270_/CLK _13271_/X VGND VGND VPWR VPWR _13254_/CLK sky130_fd_sc_hd__dlclkp_1
X_12221_ _12151_/A wr VGND VGND VPWR VPWR _12221_/X sky130_fd_sc_hd__and2_1
XFILLER_135_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[13\].VALID\[6\].TOBUF OVHB\[13\].VALID\[6\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_108_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12152_ _12151_/A VGND VGND VPWR VPWR _12152_/Y sky130_fd_sc_hd__inv_2
XOVHB\[17\].VALID\[3\].FF OVHB\[17\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[17\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11103_ _11111_/CLK line[0] VGND VGND VPWR VPWR _11103_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11809__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10713__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12109_/CLK line[64] VGND VGND VPWR VPWR _12084_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07294__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05807__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11034_ _11033_/Q _11067_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[4\].INV _13987_/X VGND VGND VPWR VPWR OVHB\[4\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[24\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12985_ _12985_/A _12992_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DEC.DEC0.AND0_A A[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11936_ _11934_/CLK line[120] VGND VGND VPWR VPWR _11936_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05542__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11867_ _11866_/Q _11872_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XMUX.MUX\[4\] _10844_/Z _05594_/Z _13504_/Z _06854_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[4] sky130_fd_sc_hd__mux4_1
X_13606_ _13598_/CLK line[115] VGND VGND VPWR VPWR _13606_/Q sky130_fd_sc_hd__dfxtp_1
X_10818_ _10804_/CLK line[121] VGND VGND VPWR VPWR _10818_/Q sky130_fd_sc_hd__dfxtp_1
X_11798_ _11776_/CLK line[57] VGND VGND VPWR VPWR _11799_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07112__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12375__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13537_ _13537_/A _13552_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_10749_ _10748_/Q _10752_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07469__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06373__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13468_ _13468_/CLK line[52] VGND VGND VPWR VPWR _13468_/Q sky130_fd_sc_hd__dfxtp_1
X_12419_ _12418_/Q _12432_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13399_ _13398_/Q _13412_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09684__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10623__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07960_ _07960_/A _07987_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09981__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05717__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06911_ _06923_/CLK line[13] VGND VGND VPWR VPWR _06911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07891_ _07905_/CLK line[77] VGND VGND VPWR VPWR _07891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09630_ _09630_/CLK _09631_/X VGND VGND VPWR VPWR _09626_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_96_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06842_ _06842_/A _06867_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07932__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[5\].FF OVHB\[15\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[15\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09561_ _09632_/A wr VGND VGND VPWR VPWR _09561_/X sky130_fd_sc_hd__and2_1
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06773_ _06775_/CLK line[78] VGND VGND VPWR VPWR _06773_/Q sky130_fd_sc_hd__dfxtp_1
X_05724_ _05724_/A _05747_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_08512_ _13921_/X VGND VGND VPWR VPWR _08512_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06548__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07006__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09492_ _09632_/A VGND VGND VPWR VPWR _09492_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[14\].FF OVHB\[31\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[31\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08443_ _08473_/CLK line[64] VGND VGND VPWR VPWR _08443_/Q sky130_fd_sc_hd__dfxtp_1
X_05655_ _05671_/CLK line[79] VGND VGND VPWR VPWR _05655_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08374_ _08373_/Q _08407_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05586_ _05586_/A _05607_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07325_ _07327_/CLK line[74] VGND VGND VPWR VPWR _07325_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13959__A A_h[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06283__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07256_ _07255_/Q _07287_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06207_ _06223_/CLK line[75] VGND VGND VPWR VPWR _06207_/Q sky130_fd_sc_hd__dfxtp_1
X_07187_ _07183_/CLK line[11] VGND VGND VPWR VPWR _07187_/Q sky130_fd_sc_hd__dfxtp_1
X_06138_ _06137_/Q _06167_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06069_ _06077_/CLK line[12] VGND VGND VPWR VPWR _06069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09828_ _09834_/CLK line[52] VGND VGND VPWR VPWR _09829_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[11\].TOBUF OVHB\[13\].VALID\[11\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_09759_ _09759_/A _09772_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11364__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11942__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06458__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12770_ _12774_/CLK line[117] VGND VGND VPWR VPWR _12770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11661__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11721_ _11720_/Q _11732_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11636_/CLK line[118] VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[7\].FF OVHB\[13\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[13\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[30\]_A3 _13599_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10603_ _10602_/Q _10612_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _11582_/Q _11592_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13308_/CLK line[113] VGND VGND VPWR VPWR _13322_/Q sky130_fd_sc_hd__dfxtp_1
X_10534_ _10520_/CLK line[119] VGND VGND VPWR VPWR _10535_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[0\].TOBUF OVHB\[28\].VALID\[0\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12923__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10465_ _10465_/A _10472_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_13253_ _13252_/Q _13272_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_12204_ _12204_/CLK line[114] VGND VGND VPWR VPWR _12204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06921__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13184_ _13194_/CLK line[50] VGND VGND VPWR VPWR _13184_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _13865_/CLK sky130_fd_sc_hd__clkbuf_4
X_10396_ _10384_/CLK line[56] VGND VGND VPWR VPWR _10396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11539__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12135_ _12134_/Q _12152_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VOBUF OVHB\[22\].V/Q OVHB\[22\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__09009__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12066_ _12072_/CLK line[51] VGND VGND VPWR VPWR _12066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11836__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13754__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11017_ _11016_/Q _11032_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08848__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12968_ _12962_/CLK line[94] VGND VGND VPWR VPWR _12969_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05272__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11919_ _11919_/A _11942_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
X_12899_ _12898_/Q _12922_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
X_05440_ _05439_/Q _05467_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08583__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05371_ _05391_/CLK line[77] VGND VGND VPWR VPWR _05371_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07199__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07110_ _07110_/CLK _07111_/X VGND VGND VPWR VPWR _07098_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07777__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08090_ _08090_/CLK _08091_/X VGND VGND VPWR VPWR _08070_/CLK sky130_fd_sc_hd__dlclkp_1
X_07041_ _07111_/A wr VGND VGND VPWR VPWR _07041_/X sky130_fd_sc_hd__and2_1
XANTENNA__07496__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[9\].FF OVHB\[11\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[11\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10353__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08992_ _08972_/CLK line[54] VGND VGND VPWR VPWR _08993_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05447__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07943_ _07942_/Q _07952_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13664__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _13480_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08758__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07874_ _07854_/CLK line[55] VGND VGND VPWR VPWR _07875_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07662__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09613_ _09612_/Q _09632_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06825_ _06825_/A _06832_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09544_ _09554_/CLK line[50] VGND VGND VPWR VPWR _09544_/Q sky130_fd_sc_hd__dfxtp_1
X_06756_ _06740_/CLK line[56] VGND VGND VPWR VPWR _06756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[3\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05707_ _05707_/A _05712_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06687_ _06687_/A _06692_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_09475_ _09474_/Q _09492_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09589__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ _08410_/CLK line[51] VGND VGND VPWR VPWR _08426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05638_ _05632_/CLK line[57] VGND VGND VPWR VPWR _05639_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05910__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10528__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ _08356_/Q _08372_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_05569_ _05568_/Q _05572_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
X_07308_ _07292_/CLK line[52] VGND VGND VPWR VPWR _07309_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08288_ _08282_/CLK line[116] VGND VGND VPWR VPWR _08288_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13839__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12743__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13201__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07239_ _07238_/Q _07252_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07837__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10250_ _10248_/CLK line[117] VGND VGND VPWR VPWR _10250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[28\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _10820_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10263__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10181_ _10180_/Q _10192_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[15\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13940_ _13944_/C _13946_/B _13944_/B _13944_/D VGND VGND VPWR VPWR _13940_/X sky130_fd_sc_hd__and4bb_4
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07572__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[1\].VALID\[2\].TOBUF OVHB\[1\].VALID\[2\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_13871_ _13870_/Q _13902_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11094__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06188__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12822_ _12820_/CLK line[27] VGND VGND VPWR VPWR _12822_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _13095_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[26\].VALID\[5\].TOBUF OVHB\[26\].VALID\[5\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09142__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12918__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12753_ _12752_/Q _12782_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09499__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11706_/CLK line[28] VGND VGND VPWR VPWR _11704_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12708_/CLK line[92] VGND VGND VPWR VPWR _12684_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05820__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[6\].VALID\[0\].FF OVHB\[6\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[6\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11635_ _11634_/Q _11662_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10438__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[17\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _11588_/CLK line[93] VGND VGND VPWR VPWR _11566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _13305_/CLK _13306_/X VGND VGND VPWR VPWR _13285_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12653__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10517_ _10517_/A _10542_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_11497_ _11497_/A _11522_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07747__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06651__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13236_ _13272_/A wr VGND VGND VPWR VPWR _13236_/X sky130_fd_sc_hd__and2_1
X_10448_ _10466_/CLK line[94] VGND VGND VPWR VPWR _10448_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11269__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ _13272_/A VGND VGND VPWR VPWR _13167_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10751__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10379_ _10379_/A _10402_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09962__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[29\].CGAND _11032_/A wr VGND VGND VPWR VPWR OVHB\[29\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09317__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12118_ _12130_/CLK line[80] VGND VGND VPWR VPWR _12118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13098_ _13120_/CLK line[16] VGND VGND VPWR VPWR _13098_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[27\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _10435_/CLK sky130_fd_sc_hd__clkbuf_4
X_04940_ A_h[9] _04940_/B2 A_h[9] _04940_/B2 VGND VGND VPWR VPWR _04940_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__10901__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12049_ _12048_/Q _12082_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08578__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09036__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06610_ _06596_/CLK line[117] VGND VGND VPWR VPWR _06611_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06098__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07590_ _07572_/CLK line[53] VGND VGND VPWR VPWR _07590_/Q sky130_fd_sc_hd__dfxtp_1
X_06541_ _06541_/A _06552_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12828__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04940__B1 A_h[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06826__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06472_ _06464_/CLK line[54] VGND VGND VPWR VPWR _06472_/Q sky130_fd_sc_hd__dfxtp_1
X_09260_ _09256_/CLK line[63] VGND VGND VPWR VPWR _09260_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09202__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08211_ _08210_/Q _08232_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_05423_ _05423_/A _05432_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_09191_ _09190_/Q _09212_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10926__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08142_ _08134_/CLK line[49] VGND VGND VPWR VPWR _08143_/A sky130_fd_sc_hd__dfxtp_1
X_05354_ _05332_/CLK line[55] VGND VGND VPWR VPWR _05354_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04924__A _04924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08073_ _08072_/Q _08092_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05285_ _05284_/Q _05292_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_07024_ _07030_/CLK line[50] VGND VGND VPWR VPWR _07024_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06561__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11179__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[2\].FF OVHB\[4\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[4\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10083__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05177__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08975_ _08974_/Q _09002_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13394__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[20\]_A2 _06539_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08488__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07926_ _07946_/CLK line[93] VGND VGND VPWR VPWR _07926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13691__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07857_ _07856_/Q _07882_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06808_ _06802_/CLK line[94] VGND VGND VPWR VPWR _06808_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[26\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _10050_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06586__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07788_ _07788_/CLK line[30] VGND VGND VPWR VPWR _07788_/Q sky130_fd_sc_hd__dfxtp_1
X_09527_ _09632_/A VGND VGND VPWR VPWR _09527_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06739_ _06738_/Q _06762_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11642__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[16\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _07180_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06736__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ _09482_/CLK line[16] VGND VGND VPWR VPWR _09458_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__04938__A1_N A_h[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09112__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08409_ _08408_/Q _08442_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10258__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XMUX.MUX\[22\] _10883_/Z _13473_/Z _06543_/Z _13613_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[22] sky130_fd_sc_hd__mux4_1
XFILLER_138_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ _09388_/Q _09422_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11420_ _11440_/CLK line[26] VGND VGND VPWR VPWR _11420_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08951__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13569__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11351_ _11351_/A _11382_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_10302_ _10314_/CLK line[27] VGND VGND VPWR VPWR _10302_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13866__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11282_ _11302_/CLK line[91] VGND VGND VPWR VPWR _11283_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13021_ _12999_/CLK line[104] VGND VGND VPWR VPWR _13021_/Q sky130_fd_sc_hd__dfxtp_1
X_10233_ _10232_/Q _10262_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05087__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].CGAND _11592_/A wr VGND VGND VPWR VPWR OVHB\[30\].CGAND/X sky130_fd_sc_hd__and2_4
X_10164_ _10188_/CLK line[92] VGND VGND VPWR VPWR _10164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11817__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10095_ _10095_/A _10122_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_13923_ _13922_/B _13923_/B _13923_/C _13923_/D VGND VGND VPWR VPWR _13923_/X sky130_fd_sc_hd__and4b_4
XOVHB\[2\].VALID\[4\].FF OVHB\[2\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[2\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ _13854_/A _13867_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12805_ _12803_/CLK line[5] VGND VGND VPWR VPWR _12805_/Q sky130_fd_sc_hd__dfxtp_1
X_13785_ _13763_/CLK line[69] VGND VGND VPWR VPWR _13785_/Q sky130_fd_sc_hd__dfxtp_1
X_10997_ _11032_/A VGND VGND VPWR VPWR _10997_/Y sky130_fd_sc_hd__inv_2
X_12736_ _12735_/Q _12747_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05550__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10168__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12667_/CLK line[70] VGND VGND VPWR VPWR _12667_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _11618_/A _11627_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[15\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _06795_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_128_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12598_ _12597_/Q _12607_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12383__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11549_ _11535_/CLK line[71] VGND VGND VPWR VPWR _11549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07477__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05070_ _05058_/CLK line[53] VGND VGND VPWR VPWR _05070_/Q sky130_fd_sc_hd__dfxtp_1
X_13219_ _13213_/CLK line[66] VGND VGND VPWR VPWR _13219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09692__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10631__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08760_ _08762_/CLK line[90] VGND VGND VPWR VPWR _08760_/Q sky130_fd_sc_hd__dfxtp_1
X_05972_ _05984_/CLK line[81] VGND VGND VPWR VPWR _05972_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[13\].TOBUF OVHB\[3\].VALID\[13\].FF/Q OVHB\[3\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05725__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08101__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07711_ _07710_/Q _07742_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_04923_ _04922_/Y _04923_/B VGND VGND VPWR VPWR _04923_/X sky130_fd_sc_hd__and2_4
X_08691_ _08690_/Q _08722_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[30\].VALID\[9\].TOBUF OVHB\[30\].VALID\[9\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_07642_ _07644_/CLK line[91] VGND VGND VPWR VPWR _07642_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07940__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[2\].TOBUF OVHB\[8\].VALID\[2\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12558__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07573_ _07572_/Q _07602_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09312_ _09311_/Q _09317_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_06524_ _06528_/CLK line[92] VGND VGND VPWR VPWR _06524_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[6\].FF OVHB\[0\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[0\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[8\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09243_ _09241_/CLK line[41] VGND VGND VPWR VPWR _09244_/A sky130_fd_sc_hd__dfxtp_1
X_06455_ _06454_/Q _06482_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09867__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05406_ _05424_/CLK line[93] VGND VGND VPWR VPWR _05406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09174_ _09173_/Q _09177_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_06386_ _06408_/CLK line[29] VGND VGND VPWR VPWR _06386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08126__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08125_ _08125_/CLK _08126_/X VGND VGND VPWR VPWR _08113_/CLK sky130_fd_sc_hd__dlclkp_1
X_05337_ _05336_/Q _05362_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12293__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10806__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06291__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[11\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08056_ _13940_/X wr VGND VGND VPWR VPWR _08056_/X sky130_fd_sc_hd__and2_1
X_05268_ _05278_/CLK line[30] VGND VGND VPWR VPWR _05268_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[14\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _06410_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11487__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07007_ _07111_/A VGND VGND VPWR VPWR _07007_/Y sky130_fd_sc_hd__inv_2
X_05199_ _05198_/Q _05222_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[7\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08958_ _08958_/A _08967_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07909_ _07905_/CLK line[71] VGND VGND VPWR VPWR _07909_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[28\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08889_ _08869_/CLK line[7] VGND VGND VPWR VPWR _08889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10920_ _10919_/Q _10927_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07850__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12468__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10851_ _10843_/CLK line[8] VGND VGND VPWR VPWR _10851_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11372__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06466__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13569_/Q _13587_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10782_ _10781_/Q _10787_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12523_/CLK line[3] VGND VGND VPWR VPWR _12521_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09777__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08681__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12452_/A _12467_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13299__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11403_ _11395_/CLK line[4] VGND VGND VPWR VPWR _11404_/A sky130_fd_sc_hd__dfxtp_1
X_12383_ _12387_/CLK line[68] VGND VGND VPWR VPWR _12383_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12781__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11334_ _11333_/Q _11347_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12931__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11265_ _11251_/CLK line[69] VGND VGND VPWR VPWR _11265_/Q sky130_fd_sc_hd__dfxtp_1
X_13004_ _13003_/Q _13027_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_10216_ _10215_/Q _10227_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_11196_ _11195_/Q _11207_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11547__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10147_ _10145_/CLK line[70] VGND VGND VPWR VPWR _10148_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09017__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[20\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10078_ _10077_/Q _10087_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08856__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _13909_/C _13909_/B _13905_/X _13909_/D VGND VGND VPWR VPWR _13552_/A sky130_fd_sc_hd__nor4b_4
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[1\].FF OVHB\[27\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[27\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13837_ _13845_/CLK line[107] VGND VGND VPWR VPWR _13837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12956__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11282__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[2\]_A2 _06780_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13768_ _13767_/Q _13797_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05280__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12719_ _12741_/CLK line[108] VGND VGND VPWR VPWR _12720_/A sky130_fd_sc_hd__dfxtp_1
X_13699_ _13701_/CLK line[44] VGND VGND VPWR VPWR _13699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06240_ _06244_/CLK line[90] VGND VGND VPWR VPWR _06240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[10\]_A1 _05576_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08591__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[30\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[24\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06171_ _06170_/Q _06202_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05122_ _05122_/CLK line[91] VGND VGND VPWR VPWR _05122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09930_ _09929_/Q _09947_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
X_05053_ _05052_/Q _05082_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[7\].TOBUF OVHB\[6\].VALID\[7\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_125_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09861_ _09849_/CLK line[67] VGND VGND VPWR VPWR _09861_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11457__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10361__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08812_ _08812_/A _08827_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_09792_ _09791_/Q _09807_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05455__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08743_ _08749_/CLK line[68] VGND VGND VPWR VPWR _08743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05955_ _05955_/CLK _05956_/X VGND VGND VPWR VPWR _05929_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[13\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13672__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13027__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08766__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08674_ _08674_/A _08687_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05886_ _13910_/X wr VGND VGND VPWR VPWR _05886_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[12\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07625_ _07633_/CLK line[69] VGND VGND VPWR VPWR _07625_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12288__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ _07555_/Q _07567_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05190__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06507_ _06489_/CLK line[70] VGND VGND VPWR VPWR _06507_/Q sky130_fd_sc_hd__dfxtp_1
X_07487_ _07467_/CLK line[6] VGND VGND VPWR VPWR _07487_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11920__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09226_ _09225_/Q _09247_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_06438_ _06437_/Q _06447_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[3\].FF OVHB\[25\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[25\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09157_ _09147_/CLK line[1] VGND VGND VPWR VPWR _09157_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10536__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06369_ _06353_/CLK line[7] VGND VGND VPWR VPWR _06369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[22\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08108_ _08108_/A _08127_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08006__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09088_ _09087_/Q _09107_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13847__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08039_ _08033_/CLK line[2] VGND VGND VPWR VPWR _08039_/Q sky130_fd_sc_hd__dfxtp_1
X_11050_ _11050_/A _11067_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10001_ _10011_/CLK line[3] VGND VGND VPWR VPWR _10001_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10271__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05365__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[5\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[11\].CGAND_A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ _11951_/Q _11977_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07580__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[2\].TOBUF OVHB\[13\].VALID\[2\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ _10903_/CLK line[46] VGND VGND VPWR VPWR _10903_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12198__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11883_ _11901_/CLK line[110] VGND VGND VPWR VPWR _11883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06196__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13622_ _13552_/A VGND VGND VPWR VPWR _13622_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10834_ _10833_/Q _10857_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13553_ _13559_/CLK line[96] VGND VGND VPWR VPWR _13553_/Q sky130_fd_sc_hd__dfxtp_1
X_10765_ _10783_/CLK line[111] VGND VGND VPWR VPWR _10765_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10296__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[14\].FF OVHB\[22\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[22\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12504_ _12503_/Q _12537_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_13484_ _13483_/Q _13517_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_10696_ _10695_/Q _10717_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_12435_ _12449_/CLK line[106] VGND VGND VPWR VPWR _12435_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10446__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12366_ _12365_/Q _12397_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_11317_ _11343_/CLK line[107] VGND VGND VPWR VPWR _11317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12661__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12297_ _12311_/CLK line[43] VGND VGND VPWR VPWR _12298_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[5\].FF OVHB\[23\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[23\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07755__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11248_ _11247_/Q _11277_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11179_ _11191_/CLK line[44] VGND VGND VPWR VPWR _11180_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09970__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05740_ _05740_/A _05747_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05671_ _05671_/CLK line[72] VGND VGND VPWR VPWR _05671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07410_ _07410_/A _07427_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
X_08390_ _08389_/Q _08407_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_07341_ _07327_/CLK line[67] VGND VGND VPWR VPWR _07341_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VOBUF OVHB\[17\].V/Q OVHB\[17\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__12836__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07272_ _07271_/Q _07287_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_09011_ _09005_/CLK line[77] VGND VGND VPWR VPWR _09011_/Q sky130_fd_sc_hd__dfxtp_1
X_06223_ _06223_/CLK line[68] VGND VGND VPWR VPWR _06223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[18\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06154_ _06154_/A _06167_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_05105_ _05093_/CLK line[69] VGND VGND VPWR VPWR _05105_/Q sky130_fd_sc_hd__dfxtp_1
X_06085_ _06077_/CLK line[5] VGND VGND VPWR VPWR _06086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09913_ _09925_/CLK line[96] VGND VGND VPWR VPWR _09913_/Q sky130_fd_sc_hd__dfxtp_1
X_05036_ _05035_/Q _05047_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11187__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09844_ _09843_/Q _09877_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09880__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09775_ _09793_/CLK line[42] VGND VGND VPWR VPWR _09775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06987_ _07001_/CLK line[33] VGND VGND VPWR VPWR _06987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13980__A A_h[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[7\].FF OVHB\[21\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[21\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08726_ _08725_/Q _08757_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08496__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05938_ _05937_/Q _05957_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[27\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08657_ _08663_/CLK line[43] VGND VGND VPWR VPWR _08657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05869_ _05871_/CLK line[34] VGND VGND VPWR VPWR _05869_/Q sky130_fd_sc_hd__dfxtp_1
X_07608_ _07608_/A _07637_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _08587_/Q _08617_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[11\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07539_ _07539_/CLK line[44] VGND VGND VPWR VPWR _07539_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11650__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].CG clk OVHB\[28\].CGAND/X VGND VGND VPWR VPWR OVHB\[28\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06744__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10550_ _10549_/Q _10577_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09120__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09209_ _09209_/A _09212_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
X_10481_ _10473_/CLK line[109] VGND VGND VPWR VPWR _10481_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _12710_/CLK sky130_fd_sc_hd__clkbuf_4
X_12220_ _12220_/CLK _12221_/X VGND VGND VPWR VPWR _12204_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13577__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[11\].VALID\[7\].TOBUF OVHB\[11\].VALID\[7\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_29_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12151_ _12151_/A wr VGND VGND VPWR VPWR _12151_/X sky130_fd_sc_hd__and2_1
X_11102_ _11032_/A VGND VGND VPWR VPWR _11102_/Y sky130_fd_sc_hd__inv_2
X_12082_ _12151_/A VGND VGND VPWR VPWR _12082_/Y sky130_fd_sc_hd__inv_2
X_11033_ _11063_/CLK line[96] VGND VGND VPWR VPWR _11033_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05095__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11825__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06919__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ _12962_/CLK line[87] VGND VGND VPWR VPWR _12985_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DEC.DEC0.AND0_B A[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11935_ _11934_/Q _11942_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11866_ _11846_/CLK line[88] VGND VGND VPWR VPWR _11866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[19\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ _13604_/Q _13622_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_10817_ _10816_/Q _10822_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11797_ _11796_/Q _11802_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11560__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13536_ _13528_/CLK line[83] VGND VGND VPWR VPWR _13537_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10748_ _10728_/CLK line[89] VGND VGND VPWR VPWR _10748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10176__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13467_ _13466_/Q _13482_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_10679_ _10678_/Q _10682_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12418_ _12414_/CLK line[84] VGND VGND VPWR VPWR _12418_/Q sky130_fd_sc_hd__dfxtp_1
X_13398_ _13394_/CLK line[20] VGND VGND VPWR VPWR _13398_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13487__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12391__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12349_ _12348_/Q _12362_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07485__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[4\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _12325_/CLK sky130_fd_sc_hd__clkbuf_4
X_06910_ _06909_/Q _06937_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_07890_ _07889_/Q _07917_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06841_ _06839_/CLK line[109] VGND VGND VPWR VPWR _06842_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11735__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[13\].TOBUF OVHB\[16\].VALID\[13\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_09560_ _09560_/CLK _09561_/X VGND VGND VPWR VPWR _09554_/CLK sky130_fd_sc_hd__dlclkp_1
X_06772_ _06771_/Q _06797_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05733__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08511_ _13921_/X wr VGND VGND VPWR VPWR _08511_/X sky130_fd_sc_hd__and2_1
X_05723_ _05739_/CLK line[110] VGND VGND VPWR VPWR _05724_/A sky130_fd_sc_hd__dfxtp_1
X_09491_ _09632_/A wr VGND VGND VPWR VPWR _09491_/X sky130_fd_sc_hd__and2_1
XFILLER_24_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08442_ _13921_/X VGND VGND VPWR VPWR _08442_/Y sky130_fd_sc_hd__inv_2
X_05654_ _05653_/Q _05677_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04927__A _04927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12566__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08373_ _08383_/CLK line[32] VGND VGND VPWR VPWR _08373_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05585_ _05575_/CLK line[47] VGND VGND VPWR VPWR _05586_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07324_ _07323_/Q _07357_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_07255_ _07267_/CLK line[42] VGND VGND VPWR VPWR _07255_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _09665_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_118_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06206_ _06205_/Q _06237_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_07186_ _07185_/Q _07217_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_06137_ _06147_/CLK line[43] VGND VGND VPWR VPWR _06137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10814__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07395__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05908__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06068_ _06067_/Q _06097_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_MUX.MUX\[23\]_A0 _13405_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05019_ _05041_/CLK line[44] VGND VGND VPWR VPWR _05019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09827_ _09827_/A _09842_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09758_ _09760_/CLK line[20] VGND VGND VPWR VPWR _09759_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05643__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08709_ _08708_/Q _08722_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_09689_ _09689_/A _09702_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[25\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11720_ _11706_/CLK line[21] VGND VGND VPWR VPWR _11720_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11651_ _11650_/Q _11662_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _10594_/CLK line[22] VGND VGND VPWR VPWR _10602_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06474__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _11588_/CLK line[86] VGND VGND VPWR VPWR _11582_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13321_ _13321_/A _13342_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10533_ _10533_/A _10542_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09785__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13252_ _13254_/CLK line[81] VGND VGND VPWR VPWR _13252_/Q sky130_fd_sc_hd__dfxtp_1
X_10464_ _10466_/CLK line[87] VGND VGND VPWR VPWR _10465_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12203_ _12202_/Q _12222_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[1\].TOBUF OVHB\[26\].VALID\[1\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10724__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13183_ _13182_/Q _13202_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_10395_ _10394_/Q _10402_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13100__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05818__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12134_ _12130_/CLK line[82] VGND VGND VPWR VPWR _12134_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _09280_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_78_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12065_ _12064_/Q _12082_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11016_ _11002_/CLK line[83] VGND VGND VPWR VPWR _11016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06649__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09025__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12967_ _12967_/A _12992_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11918_ _11934_/CLK line[126] VGND VGND VPWR VPWR _11919_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12898_ _12902_/CLK line[62] VGND VGND VPWR VPWR _12898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11849_ _11848_/Q _11872_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11290__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].CGAND _09912_/A wr VGND VGND VPWR VPWR OVHB\[25\].CG/GATE sky130_fd_sc_hd__and2_4
XFILLER_53_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06384__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05370_ _05369_/Q _05397_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_13519_ _13518_/Q _13552_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07040_ _07040_/CLK _07041_/X VGND VGND VPWR VPWR _07030_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_115_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08991_ _08991_/A _09002_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[18\].VALID\[7\].TOBUF OVHB\[18\].VALID\[7\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_07942_ _07946_/CLK line[86] VGND VGND VPWR VPWR _07942_/Q sky130_fd_sc_hd__dfxtp_1
X_07873_ _07872_/Q _07882_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06202__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11465__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[7\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[22\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _08895_/CLK sky130_fd_sc_hd__clkbuf_4
X_09612_ _09626_/CLK line[81] VGND VGND VPWR VPWR _09612_/Q sky130_fd_sc_hd__dfxtp_1
X_06824_ _06802_/CLK line[87] VGND VGND VPWR VPWR _06825_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06559__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05463__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[12\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _06025_/CLK sky130_fd_sc_hd__clkbuf_4
X_09543_ _09542_/Q _09562_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_06755_ _06754_/Q _06762_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13680__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05706_ _05708_/CLK line[88] VGND VGND VPWR VPWR _05707_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08774__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09474_ _09482_/CLK line[18] VGND VGND VPWR VPWR _09474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06686_ _06682_/CLK line[24] VGND VGND VPWR VPWR _06687_/A sky130_fd_sc_hd__dfxtp_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ _08425_/A _08442_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_05637_ _05637_/A _05642_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _08358_/CLK line[19] VGND VGND VPWR VPWR _08356_/Q sky130_fd_sc_hd__dfxtp_1
X_05568_ _05568_/CLK line[25] VGND VGND VPWR VPWR _05568_/Q sky130_fd_sc_hd__dfxtp_1
X_07307_ _07306_/Q _07322_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_08287_ _08286_/Q _08302_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_05499_ _05498_/Q _05502_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_07238_ _07232_/CLK line[20] VGND VGND VPWR VPWR _07238_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].INV _13986_/X VGND VGND VPWR VPWR OVHB\[3\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_118_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07169_ _07168_/Q _07182_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05638__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08014__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10180_ _10188_/CLK line[85] VGND VGND VPWR VPWR _10180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13855__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08949__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13870_ _13882_/CLK line[122] VGND VGND VPWR VPWR _13870_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05373__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[14\].FF OVHB\[27\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[27\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12821_ _12821_/A _12852_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13590__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[24\].VALID\[6\].TOBUF OVHB\[24\].VALID\[6\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12752_ _12774_/CLK line[123] VGND VGND VPWR VPWR _12752_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11702_/Q _11732_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12682_/Q _12712_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _05640_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11636_/CLK line[124] VGND VGND VPWR VPWR _11634_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[23\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _11564_/Q _11592_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13304_ _13303_/Q _13307_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10516_ _10520_/CLK line[125] VGND VGND VPWR VPWR _10517_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11496_ _11500_/CLK line[61] VGND VGND VPWR VPWR _11497_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13235_ _13235_/CLK _13236_/X VGND VGND VPWR VPWR _13213_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10454__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[5\].FF OVHB\[9\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[9\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10447_ _10446_/Q _10472_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05548__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13166_ _13272_/A wr VGND VGND VPWR VPWR _13166_/X sky130_fd_sc_hd__and2_1
X_10378_ _10384_/CLK line[62] VGND VGND VPWR VPWR _10379_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13765__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10751__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12117_ _12151_/A VGND VGND VPWR VPWR _12117_/Y sky130_fd_sc_hd__inv_2
X_13097_ _13272_/A VGND VGND VPWR VPWR _13097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07763__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12048_ _12072_/CLK line[48] VGND VGND VPWR VPWR _12048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[5\]_A0 _10846_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06540_ _06528_/CLK line[85] VGND VGND VPWR VPWR _06541_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04940__B2 _04940_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06471_ _06470_/Q _06482_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10629__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13005__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08210_ _08208_/CLK line[95] VGND VGND VPWR VPWR _08210_/Q sky130_fd_sc_hd__dfxtp_1
X_05422_ _05424_/CLK line[86] VGND VGND VPWR VPWR _05423_/A sky130_fd_sc_hd__dfxtp_1
X_09190_ _09200_/CLK line[31] VGND VGND VPWR VPWR _09190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06692__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07003__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10926__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].V OVHB\[6\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[6\].V/Q sky130_fd_sc_hd__dfrtp_1
X_08141_ _08140_/Q _08162_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_05353_ _05352_/Q _05362_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12844__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07938__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[10\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _05255_/CLK sky130_fd_sc_hd__clkbuf_4
X_08072_ _08070_/CLK line[17] VGND VGND VPWR VPWR _08072_/Q sky130_fd_sc_hd__dfxtp_1
X_05284_ _05278_/CLK line[23] VGND VGND VPWR VPWR _05284_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[5\].TOBUF OVHB\[30\].VALID\[5\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_07023_ _07022_/Q _07042_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08974_ _08972_/CLK line[60] VGND VGND VPWR VPWR _08974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[6\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07673__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[20\]_A3 _07169_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07925_ _07924_/Q _07952_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11195__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[7\].VALID\[7\].FF OVHB\[7\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[7\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06289__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07856_ _07854_/CLK line[61] VGND VGND VPWR VPWR _07856_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06867__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06807_ _06806_/Q _06832_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07787_ _07786_/Q _07812_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06586__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04999_ _04998_/Q _05012_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_09526_ _09632_/A wr VGND VGND VPWR VPWR _09526_/X sky130_fd_sc_hd__and2_1
X_06738_ _06740_/CLK line[62] VGND VGND VPWR VPWR _06738_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09457_ _09632_/A VGND VGND VPWR VPWR _09457_/Y sky130_fd_sc_hd__inv_2
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06669_ _06668_/Q _06692_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08408_ _08410_/CLK line[48] VGND VGND VPWR VPWR _08408_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09388_ _09414_/CLK line[112] VGND VGND VPWR VPWR _09388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XMUX.MUX\[15\] _11396_/Z _05586_/Z _13496_/Z _13566_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[15] sky130_fd_sc_hd__mux4_1
XANTENNA__12754__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08339_ _08338_/Q _08372_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07848__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06752__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11350_ _11370_/CLK line[122] VGND VGND VPWR VPWR _11351_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05011__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10301_ _10300_/Q _10332_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_11281_ _11280_/Q _11312_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13020_ _13019_/Q _13027_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_10232_ _10248_/CLK line[123] VGND VGND VPWR VPWR _10232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08679__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10163_ _10163_/A _10192_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10094_ _10100_/CLK line[60] VGND VGND VPWR VPWR _10095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13922_ _13923_/B _13922_/B _13923_/C _13923_/D VGND VGND VPWR VPWR _13922_/X sky130_fd_sc_hd__and4b_4
XANTENNA_OVHB\[12\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].V OVHB\[20\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[20\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ _13845_/CLK line[100] VGND VGND VPWR VPWR _13854_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12929__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11833__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12804_ _12804_/A _12817_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06927__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13784_ _13783_/Q _13797_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10996_ _11032_/A wr VGND VGND VPWR VPWR _10996_/X sky130_fd_sc_hd__and2_1
XANTENNA__09303__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[9\].FF OVHB\[5\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[5\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12735_ _12741_/CLK line[101] VGND VGND VPWR VPWR _12735_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12665_/Q _12677_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _11605_/CLK line[102] VGND VGND VPWR VPWR _11618_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12601_/CLK line[38] VGND VGND VPWR VPWR _12597_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06662__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11548_ _11547_/Q _11557_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10184__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[11\].TOBUF OVHB\[26\].VALID\[11\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_11479_ _11479_/CLK line[39] VGND VGND VPWR VPWR _11479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05278__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13218_ _13218_/A _13237_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08232__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[21\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13495__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[23\].VALID\[12\].FF OVHB\[23\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[23\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13149_ _13163_/CLK line[34] VGND VGND VPWR VPWR _13149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08589__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07493__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05971_ _05970_/Q _05992_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_07710_ _07724_/CLK line[122] VGND VGND VPWR VPWR _07710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04922_ A_h[23] VGND VGND VPWR VPWR _04922_/Y sky130_fd_sc_hd__inv_2
X_08690_ _08710_/CLK line[58] VGND VGND VPWR VPWR _08690_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].V OVHB\[11\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[11\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07641_ _07641_/A _07672_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11743__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07572_ _07572_/CLK line[59] VGND VGND VPWR VPWR _07572_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06837__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05741__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09213__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09311_ _09307_/CLK line[72] VGND VGND VPWR VPWR _09311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06523_ _06522_/Q _06552_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[3\].TOBUF OVHB\[6\].VALID\[3\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10359__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[4\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09242_ _09242_/A _09247_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_06454_ _06464_/CLK line[60] VGND VGND VPWR VPWR _06454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08407__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05405_ _05404_/Q _05432_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_09173_ _09147_/CLK line[9] VGND VGND VPWR VPWR _09173_/Q sky130_fd_sc_hd__dfxtp_1
X_06385_ _06384_/Q _06412_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[14\].FF OVHB\[13\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[13\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08126__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07668__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08124_ _08123_/Q _08127_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_05336_ _05332_/CLK line[61] VGND VGND VPWR VPWR _05336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10094__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08055_ _08055_/CLK _08056_/X VGND VGND VPWR VPWR _08033_/CLK sky130_fd_sc_hd__dlclkp_1
X_05267_ _05266_/Q _05292_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05188__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07006_ _07111_/A wr VGND VGND VPWR VPWR _07006_/X sky130_fd_sc_hd__and2_1
X_05198_ _05214_/CLK line[126] VGND VGND VPWR VPWR _05198_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11918__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05916__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08957_ _08947_/CLK line[38] VGND VGND VPWR VPWR _08958_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07908_ _07907_/Q _07917_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
X_08888_ _08888_/A _08897_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_07839_ _07837_/CLK line[39] VGND VGND VPWR VPWR _07839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ _10850_/A _10857_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05651__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[18\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09701__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09509_ _09507_/CLK line[34] VGND VGND VPWR VPWR _09509_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10269__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10781_ _10783_/CLK line[104] VGND VGND VPWR VPWR _10781_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A _12537_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[14\].VALID\[1\].FF OVHB\[14\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[14\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12449_/CLK line[99] VGND VGND VPWR VPWR _12452_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12484__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[5\].FF OVHB\[31\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[31\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07578__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11402_ _11401_/Q _11417_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_12382_ _12381_/Q _12397_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12781__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11333_ _11343_/CLK line[100] VGND VGND VPWR VPWR _11333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09793__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05676__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11264_ _11263_/Q _11277_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13003_ _12999_/CLK line[110] VGND VGND VPWR VPWR _13003_/Q sky130_fd_sc_hd__dfxtp_1
X_10215_ _10217_/CLK line[101] VGND VGND VPWR VPWR _10215_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10732__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11195_ _11191_/CLK line[37] VGND VGND VPWR VPWR _11195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05826__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10146_ _10145_/Q _10157_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08202__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10077_ _10073_/CLK line[38] VGND VGND VPWR VPWR _10077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13905_ A[6] VGND VGND VPWR VPWR _13905_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12659__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13836_ _13836_/A _13867_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09033__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[2\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _11380_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__12956__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[2\]_A3 _13570_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _13763_/CLK line[75] VGND VGND VPWR VPWR _13767_/Q sky130_fd_sc_hd__dfxtp_1
X_10979_ _10977_/CLK line[66] VGND VGND VPWR VPWR _10979_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09968__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12718_ _12717_/Q _12747_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_13698_ _13697_/Q _13727_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10907__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[10\]_A2 _13486_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12649_ _12667_/CLK line[76] VGND VGND VPWR VPWR _12649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06392__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06170_ _06186_/CLK line[58] VGND VGND VPWR VPWR _06170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05121_ _05120_/Q _05152_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[12\].VALID\[3\].FF OVHB\[12\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[12\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05052_ _05058_/CLK line[59] VGND VGND VPWR VPWR _05052_/Q sky130_fd_sc_hd__dfxtp_1
X_09860_ _09860_/A _09877_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[4\].VALID\[8\].TOBUF OVHB\[4\].VALID\[8\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08897__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09208__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VOBUF OVHB\[13\].V/Q OVHB\[13\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_98_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08811_ _08823_/CLK line[99] VGND VGND VPWR VPWR _08812_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04937__A1_N A_h[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09791_ _09793_/CLK line[35] VGND VGND VPWR VPWR _09791_/Q sky130_fd_sc_hd__dfxtp_1
X_08742_ _08741_/Q _08757_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_05954_ _05953_/Q _05957_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08673_ _08663_/CLK line[36] VGND VGND VPWR VPWR _08674_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05885_ _05885_/CLK _05886_/X VGND VGND VPWR VPWR _05871_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11473__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07624_ _07623_/Q _07637_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06567__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _07539_/CLK line[37] VGND VGND VPWR VPWR _07555_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09878__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06506_ _06505_/Q _06517_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08782__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07486_ _07486_/A _07497_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09225_ _09241_/CLK line[47] VGND VGND VPWR VPWR _09225_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07041__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06437_ _06421_/CLK line[38] VGND VGND VPWR VPWR _06437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[1\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _08195_/CLK sky130_fd_sc_hd__clkbuf_4
X_09156_ _09155_/Q _09177_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_06368_ _06368_/A _06377_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_08107_ _08113_/CLK line[33] VGND VGND VPWR VPWR _08108_/A sky130_fd_sc_hd__dfxtp_1
X_05319_ _05299_/CLK line[39] VGND VGND VPWR VPWR _05319_/Q sky130_fd_sc_hd__dfxtp_1
X_09087_ _09085_/CLK line[97] VGND VGND VPWR VPWR _09087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06299_ _06285_/CLK line[103] VGND VGND VPWR VPWR _06299_/Q sky130_fd_sc_hd__dfxtp_1
X_08038_ _08037_/Q _08057_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[8\].FF OVHB\[28\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[28\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11648__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09118__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10000_ _10000_/A _10017_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13863__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09989_ _10011_/CLK line[12] VGND VGND VPWR VPWR _09989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08957__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[5\].FF OVHB\[10\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[10\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07216__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[31\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _11765_/CLK sky130_fd_sc_hd__clkbuf_4
X_11951_ _11945_/CLK line[13] VGND VGND VPWR VPWR _11951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11383__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10902_ _10902_/A _10927_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[3\].TOBUF OVHB\[11\].VALID\[3\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_11882_ _11881_/Q _11907_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].CGAND_A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05381__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10833_ _10843_/CLK line[14] VGND VGND VPWR VPWR _10833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13621_ _13552_/A wr VGND VGND VPWR VPWR _13621_/X sky130_fd_sc_hd__and2_1
XANTENNA__10577__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08692__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _13552_/A VGND VGND VPWR VPWR _13552_/Y sky130_fd_sc_hd__inv_2
X_10764_ _10763_/Q _10787_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10296__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DECH.DEC0.AND3_A A_h[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12503_ _12523_/CLK line[0] VGND VGND VPWR VPWR _12503_/Q sky130_fd_sc_hd__dfxtp_1
X_13483_ _13497_/CLK line[64] VGND VGND VPWR VPWR _13483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10695_ _10707_/CLK line[79] VGND VGND VPWR VPWR _10695_/Q sky130_fd_sc_hd__dfxtp_1
X_12434_ _12433_/Q _12467_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12365_ _12387_/CLK line[74] VGND VGND VPWR VPWR _12365_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[0\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _05010_/CLK sky130_fd_sc_hd__clkbuf_4
X_11316_ _11315_/Q _11347_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06940__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12296_ _12295_/Q _12327_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11558__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10462__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11247_ _11251_/CLK line[75] VGND VGND VPWR VPWR _11247_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05556__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11178_ _11178_/A _11207_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13773__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10129_ _10145_/CLK line[76] VGND VGND VPWR VPWR _10129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08867__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07771__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12389__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11871__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05670_ _05670_/A _05677_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13819_ _13818_/Q _13832_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09698__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07340_ _07339_/Q _07357_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07271_ _07267_/CLK line[35] VGND VGND VPWR VPWR _07271_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10637__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[20\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _08510_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13013__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09010_ _09009_/Q _09037_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_06222_ _06221_/Q _06237_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08107__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[18\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06153_ _06147_/CLK line[36] VGND VGND VPWR VPWR _06154_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07946__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05104_ _05103_/Q _05117_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_06084_ _06083_/Q _06097_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[21\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05035_ _05041_/CLK line[37] VGND VGND VPWR VPWR _05035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10372__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09912_ _09912_/A VGND VGND VPWR VPWR _09912_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09843_ _09849_/CLK line[64] VGND VGND VPWR VPWR _09843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09774_ _09773_/Q _09807_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_06986_ _06986_/A _07007_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07681__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12299__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05937_ _05929_/CLK line[65] VGND VGND VPWR VPWR _05937_/Q sky130_fd_sc_hd__dfxtp_1
X_08725_ _08749_/CLK line[74] VGND VGND VPWR VPWR _08725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06297__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08656_ _08655_/Q _08687_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05868_ _05868_/A _05887_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07607_ _07633_/CLK line[75] VGND VGND VPWR VPWR _07608_/A sky130_fd_sc_hd__dfxtp_1
X_08587_ _08609_/CLK line[11] VGND VGND VPWR VPWR _08587_/Q sky130_fd_sc_hd__dfxtp_1
X_05799_ _05799_/CLK line[2] VGND VGND VPWR VPWR _05800_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ _07537_/Q _07567_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[4\].VALID\[14\].FF OVHB\[4\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[4\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10547__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07469_ _07467_/CLK line[12] VGND VGND VPWR VPWR _07469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ _09200_/CLK line[25] VGND VGND VPWR VPWR _09209_/A sky130_fd_sc_hd__dfxtp_1
X_10480_ _10479_/Q _10507_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_09139_ _09138_/Q _09142_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12762__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12117__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07856__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ _12150_/CLK _12151_/X VGND VGND VPWR VPWR _12130_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11378__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11101_ _11032_/A wr VGND VGND VPWR VPWR _11101_/X sky130_fd_sc_hd__and2_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12081_ _12151_/A wr VGND VGND VPWR VPWR _12081_/X sky130_fd_sc_hd__and2_1
X_11032_ _11032_/A VGND VGND VPWR VPWR _11032_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12983_ _12982_/Q _12992_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12002__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11934_ _11934_/CLK line[119] VGND VGND VPWR VPWR _11934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[2\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12937__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11865_ _11864_/Q _11872_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_13604_ _13598_/CLK line[114] VGND VGND VPWR VPWR _13604_/Q sky130_fd_sc_hd__dfxtp_1
X_10816_ _10804_/CLK line[120] VGND VGND VPWR VPWR _10816_/Q sky130_fd_sc_hd__dfxtp_1
X_11796_ _11776_/CLK line[56] VGND VGND VPWR VPWR _11796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09311__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13535_ _13535_/A _13552_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_10747_ _10746_/Q _10752_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13411__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[12\].FF OVHB\[28\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[28\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10678_ _10656_/CLK line[57] VGND VGND VPWR VPWR _10678_/Q sky130_fd_sc_hd__dfxtp_1
X_13466_ _13468_/CLK line[51] VGND VGND VPWR VPWR _13466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12417_ _12416_/Q _12432_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13397_ _13396_/Q _13412_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06670__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12348_ _12352_/CLK line[52] VGND VGND VPWR VPWR _12348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11288__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[14\].TOBUF OVHB\[12\].VALID\[14\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_12279_ _12279_/A _12292_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05286__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].CGAND _13922_/X wr VGND VGND VPWR VPWR OVHB\[21\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06840_ _06839_/Q _06867_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08597__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06771_ _06775_/CLK line[77] VGND VGND VPWR VPWR _06771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08510_ _08510_/CLK _08511_/X VGND VGND VPWR VPWR _08480_/CLK sky130_fd_sc_hd__dlclkp_1
X_05722_ _05721_/Q _05747_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_09490_ _09490_/CLK _09491_/X VGND VGND VPWR VPWR _09482_/CLK sky130_fd_sc_hd__dlclkp_1
X_08441_ _13921_/X wr VGND VGND VPWR VPWR _08441_/X sky130_fd_sc_hd__and2_1
XANTENNA__09071__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[14\].FF OVHB\[18\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[18\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05653_ _05671_/CLK line[78] VGND VGND VPWR VPWR _05653_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11751__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06845__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08372_ _13921_/X VGND VGND VPWR VPWR _08372_/Y sky130_fd_sc_hd__inv_2
X_05584_ _05583_/Q _05607_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[3\].TOBUF OVHB\[18\].VALID\[3\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__09221__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[0\].FF OVHB\[1\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[1\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07323_ _07327_/CLK line[64] VGND VGND VPWR VPWR _07323_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[12\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07254_ _07253_/Q _07287_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13678__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06205_ _06223_/CLK line[74] VGND VGND VPWR VPWR _06205_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[17\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07185_ _07183_/CLK line[10] VGND VGND VPWR VPWR _07185_/Q sky130_fd_sc_hd__dfxtp_1
X_06136_ _06136_/A _06167_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[23\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06067_ _06077_/CLK line[11] VGND VGND VPWR VPWR _06067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05196__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[23\]_A1 _09555_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09246__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05018_ _05017_/Q _05047_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11926__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09826_ _09834_/CLK line[51] VGND VGND VPWR VPWR _09827_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[5\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09757_ _09756_/Q _09772_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_06969_ _06969_/A _06972_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
X_08708_ _08710_/CLK line[52] VGND VGND VPWR VPWR _08708_/Q sky130_fd_sc_hd__dfxtp_1
X_09688_ _09694_/CLK line[116] VGND VGND VPWR VPWR _09689_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[31\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08639_ _08638_/Q _08652_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11636_/CLK line[117] VGND VGND VPWR VPWR _11650_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[8\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10277__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _10600_/Q _10612_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _11580_/Q _11592_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08970__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13308_/CLK line[127] VGND VGND VPWR VPWR _13321_/A sky130_fd_sc_hd__dfxtp_1
X_10532_ _10520_/CLK line[118] VGND VGND VPWR VPWR _10533_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13588__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12492__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10463_ _10462_/Q _10472_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_13251_ _13250_/Q _13272_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07586__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12202_ _12204_/CLK line[113] VGND VGND VPWR VPWR _12202_/Q sky130_fd_sc_hd__dfxtp_1
X_13182_ _13194_/CLK line[49] VGND VGND VPWR VPWR _13182_/Q sky130_fd_sc_hd__dfxtp_1
X_10394_ _10384_/CLK line[55] VGND VGND VPWR VPWR _10394_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[2\].TOBUF OVHB\[24\].VALID\[2\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_12133_ _12133_/A _12152_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_12064_ _12072_/CLK line[50] VGND VGND VPWR VPWR _12064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11015_ _11014_/Q _11032_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10740__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05834__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[12\].FF OVHB\[0\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[0\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08210__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12966_ _12962_/CLK line[93] VGND VGND VPWR VPWR _12967_/A sky130_fd_sc_hd__dfxtp_1
X_11917_ _11916_/Q _11942_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12667__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12897_ _12896_/Q _12922_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11848_ _11846_/CLK line[94] VGND VGND VPWR VPWR _11848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11779_ _11778_/Q _11802_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09976__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13518_ _13528_/CLK line[80] VGND VGND VPWR VPWR _13518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10915__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13449_ _13448_/Q _13482_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _08972_/CLK line[53] VGND VGND VPWR VPWR _08991_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07941_ _07941_/A _07952_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[16\].VALID\[8\].TOBUF OVHB\[16\].VALID\[8\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10650__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07872_ _07854_/CLK line[54] VGND VGND VPWR VPWR _07872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[18\].CG clk OVHB\[18\].CGAND/X VGND VGND VPWR VPWR OVHB\[18\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09611_ _09610_/Q _09632_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_06823_ _06822_/Q _06832_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[30\].VALID\[1\].TOBUF OVHB\[30\].VALID\[1\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_110_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06754_ _06740_/CLK line[55] VGND VGND VPWR VPWR _06754_/Q sky130_fd_sc_hd__dfxtp_1
X_09542_ _09554_/CLK line[49] VGND VGND VPWR VPWR _09542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05705_ _05704_/Q _05712_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12577__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[10\].FF OVHB\[24\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[24\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06685_ _06685_/A _06692_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_09473_ _09473_/A _09492_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11481__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05636_ _05632_/CLK line[56] VGND VGND VPWR VPWR _05637_/A sky130_fd_sc_hd__dfxtp_1
X_08424_ _08410_/CLK line[50] VGND VGND VPWR VPWR _08425_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06575__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _08355_/A _08372_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05567_ _05567_/A _05572_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09886__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07306_ _07292_/CLK line[51] VGND VGND VPWR VPWR _07306_/Q sky130_fd_sc_hd__dfxtp_1
X_08286_ _08282_/CLK line[115] VGND VGND VPWR VPWR _08286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05498_ _05476_/CLK line[121] VGND VGND VPWR VPWR _05498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10825__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07237_ _07236_/Q _07252_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_07168_ _07170_/CLK line[116] VGND VGND VPWR VPWR _07168_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[10\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06119_ _06118_/Q _06132_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_07099_ _07099_/A _07112_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11656__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[12\].FF OVHB\[14\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[14\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09126__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09809_ _09809_/A _09842_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12820_ _12820_/CLK line[26] VGND VGND VPWR VPWR _12821_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12750_/Q _12782_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11391__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[3\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06485__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11702_ _11706_/CLK line[27] VGND VGND VPWR VPWR _11702_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[7\].TOBUF OVHB\[22\].VALID\[7\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12708_/CLK line[91] VGND VGND VPWR VPWR _12682_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11633_ _11632_/Q _11662_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[6\].VALID\[11\].TOBUF OVHB\[6\].VALID\[11\].FF/Q OVHB\[6\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _11588_/CLK line[92] VGND VGND VPWR VPWR _11564_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13285_/CLK line[105] VGND VGND VPWR VPWR _13303_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10515_ _10514_/Q _10542_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_11495_ _11494_/Q _11522_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_13234_ _13233_/Q _13237_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_10446_ _10466_/CLK line[93] VGND VGND VPWR VPWR _10446_/Q sky130_fd_sc_hd__dfxtp_1
X_13165_ _13165_/CLK _13166_/X VGND VGND VPWR VPWR _13163_/CLK sky130_fd_sc_hd__dlclkp_1
X_10377_ _10376_/Q _10402_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12116_ _12151_/A wr VGND VGND VPWR VPWR _12116_/X sky130_fd_sc_hd__and2_1
X_13096_ _13272_/A wr VGND VGND VPWR VPWR _13096_/X sky130_fd_sc_hd__and2_1
XANTENNA__11566__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12047_ _12151_/A VGND VGND VPWR VPWR _12047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05564__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13781__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08875__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[5\]_A1 _05036_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12949_ _12937_/CLK line[71] VGND VGND VPWR VPWR _12949_/Q sky130_fd_sc_hd__dfxtp_1
X_06470_ _06464_/CLK line[53] VGND VGND VPWR VPWR _06470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[13\]_A0 _13352_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05421_ _05420_/Q _05432_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08140_ _08134_/CLK line[63] VGND VGND VPWR VPWR _08140_/Q sky130_fd_sc_hd__dfxtp_1
X_05352_ _05332_/CLK line[54] VGND VGND VPWR VPWR _05352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08071_ _08070_/Q _08092_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_05283_ _05282_/Q _05292_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13021__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05739__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07022_ _07030_/CLK line[49] VGND VGND VPWR VPWR _07022_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08115__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08973_ _08972_/Q _09002_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10380__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07924_ _07946_/CLK line[92] VGND VGND VPWR VPWR _07924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05474__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07855_ _07855_/A _07882_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[14\].FF OVHB\[9\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[9\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06806_ _06802_/CLK line[93] VGND VGND VPWR VPWR _06806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[22\].VALID\[1\].FF OVHB\[22\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[22\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07786_ _07788_/CLK line[29] VGND VGND VPWR VPWR _07786_/Q sky130_fd_sc_hd__dfxtp_1
X_04998_ _05000_/CLK line[20] VGND VGND VPWR VPWR _04998_/Q sky130_fd_sc_hd__dfxtp_1
X_09525_ _09525_/CLK _09526_/X VGND VGND VPWR VPWR _09507_/CLK sky130_fd_sc_hd__dlclkp_1
X_06737_ _06736_/Q _06762_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ _09632_/A wr VGND VGND VPWR VPWR _09456_/X sky130_fd_sc_hd__and2_1
X_06668_ _06682_/CLK line[30] VGND VGND VPWR VPWR _06668_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05619_ _05618_/Q _05642_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08407_ _13921_/X VGND VGND VPWR VPWR _08407_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09387_ _09352_/A VGND VGND VPWR VPWR _09387_/Y sky130_fd_sc_hd__inv_2
X_06599_ _06599_/A _06622_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08338_ _08358_/CLK line[16] VGND VGND VPWR VPWR _08338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10555__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08269_ _08268_/Q _08302_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05649__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10300_ _10314_/CLK line[26] VGND VGND VPWR VPWR _10300_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05011__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08025__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11280_ _11302_/CLK line[90] VGND VGND VPWR VPWR _11280_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[13\].TOBUF OVHB\[29\].VALID\[13\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_10231_ _10230_/Q _10262_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12770__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07864__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _10188_/CLK line[91] VGND VGND VPWR VPWR _10163_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10093_ _10092_/Q _10122_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13921_ _13922_/B _13923_/B _13923_/C _13923_/D VGND VGND VPWR VPWR _13921_/X sky130_fd_sc_hd__and4bb_4
X_13852_ _13852_/A _13867_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12803_ _12803_/CLK line[4] VGND VGND VPWR VPWR _12804_/A sky130_fd_sc_hd__dfxtp_1
X_13783_ _13763_/CLK line[68] VGND VGND VPWR VPWR _13783_/Q sky130_fd_sc_hd__dfxtp_1
X_10995_ _10995_/CLK _10996_/X VGND VGND VPWR VPWR _10977_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13106__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _12734_/A _12747_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07104__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12945__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[12\].TOBUF OVHB\[22\].VALID\[12\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12667_/CLK line[69] VGND VGND VPWR VPWR _12665_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[3\].FF OVHB\[20\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[20\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _11615_/Q _11627_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A _12607_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _11535_/CLK line[70] VGND VGND VPWR VPWR _11547_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[10\].VALID\[10\].FF OVHB\[10\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[10\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11478_ _11477_/Q _11487_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_13217_ _13213_/CLK line[65] VGND VGND VPWR VPWR _13218_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12680__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10429_ _10405_/CLK line[71] VGND VGND VPWR VPWR _10429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13148_ _13147_/Q _13167_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11296__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05970_ _05984_/CLK line[95] VGND VGND VPWR VPWR _05970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13079_ _13075_/CLK line[2] VGND VGND VPWR VPWR _13079_/Q sky130_fd_sc_hd__dfxtp_1
X_04921_ _04916_/X _04918_/Y _04921_/C _04921_/D VGND VGND VPWR VPWR _04921_/X sky130_fd_sc_hd__and4_4
XFILLER_39_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07640_ _07644_/CLK line[90] VGND VGND VPWR VPWR _07641_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].INV _13985_/X VGND VGND VPWR VPWR OVHB\[2\].INV/Y sky130_fd_sc_hd__inv_2
X_07571_ _07570_/Q _07602_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06522_ _06528_/CLK line[91] VGND VGND VPWR VPWR _06522_/Q sky130_fd_sc_hd__dfxtp_1
X_09310_ _09309_/Q _09317_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07014__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[4\].TOBUF OVHB\[4\].VALID\[4\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[4\].FF OVHB\[19\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[19\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06453_ _06453_/A _06482_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
X_09241_ _09241_/CLK line[40] VGND VGND VPWR VPWR _09242_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12855__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[7\].TOBUF OVHB\[29\].VALID\[7\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_05404_ _05424_/CLK line[92] VGND VGND VPWR VPWR _05404_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06853__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09172_ _09171_/Q _09177_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_06384_ _06408_/CLK line[28] VGND VGND VPWR VPWR _06384_/Q sky130_fd_sc_hd__dfxtp_1
X_08123_ _08113_/CLK line[41] VGND VGND VPWR VPWR _08123_/Q sky130_fd_sc_hd__dfxtp_1
X_05335_ _05334_/Q _05362_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ _08053_/Q _08057_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05266_ _05278_/CLK line[29] VGND VGND VPWR VPWR _05266_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13686__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07005_ _07005_/CLK _07006_/X VGND VGND VPWR VPWR _07001_/CLK sky130_fd_sc_hd__dlclkp_1
X_05197_ _05196_/Q _05222_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08956_ _08955_/Q _08967_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05782__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07907_ _07905_/CLK line[70] VGND VGND VPWR VPWR _07907_/Q sky130_fd_sc_hd__dfxtp_1
X_08887_ _08869_/CLK line[6] VGND VGND VPWR VPWR _08888_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11934__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07838_ _07838_/A _07847_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09404__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07769_ _07773_/CLK line[7] VGND VGND VPWR VPWR _07770_/A sky130_fd_sc_hd__dfxtp_1
X_09508_ _09508_/A _09527_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09701__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10780_ _10779_/Q _10787_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _09427_/CLK line[2] VGND VGND VPWR VPWR _09440_/A sky130_fd_sc_hd__dfxtp_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12449_/Q _12467_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06763__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10285__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11401_ _11395_/CLK line[3] VGND VGND VPWR VPWR _11401_/Q sky130_fd_sc_hd__dfxtp_1
X_12381_ _12387_/CLK line[67] VGND VGND VPWR VPWR _12381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05379__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05957__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11332_ _11332_/A _11347_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[17\].VALID\[6\].FF OVHB\[17\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[17\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13596__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[26\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05676__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11263_ _11251_/CLK line[68] VGND VGND VPWR VPWR _11263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[5\].VALID\[12\].FF OVHB\[5\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[5\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07594__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13002_ _13001_/Q _13027_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_10214_ _10213_/Q _10227_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_11194_ _11193_/Q _11207_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10145_ _10145_/CLK line[69] VGND VGND VPWR VPWR _10145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06003__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10076_ _10075_/Q _10087_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11844__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13904_ A[5] VGND VGND VPWR VPWR _13909_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__06938__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05842__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13835_ _13845_/CLK line[106] VGND VGND VPWR VPWR _13836_/A sky130_fd_sc_hd__dfxtp_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ _13765_/Q _13797_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_10978_ _10978_/A _10997_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_12717_ _12741_/CLK line[107] VGND VGND VPWR VPWR _12717_/Q sky130_fd_sc_hd__dfxtp_1
X_13697_ _13701_/CLK line[43] VGND VGND VPWR VPWR _13697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07769__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12648_ _12647_/Q _12677_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[10\]_A3 _07116_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10195__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12579_ _12601_/CLK line[44] VGND VGND VPWR VPWR _12580_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05120_ _05122_/CLK line[90] VGND VGND VPWR VPWR _05120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10923__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05051_ _05050_/Q _05082_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[2\].VALID\[9\].TOBUF OVHB\[2\].VALID\[9\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_08810_ _08809_/Q _08827_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09790_ _09789_/Q _09807_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[8\].FF OVHB\[15\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[15\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__04919__A2_N _04919_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[10\].FF OVHB\[29\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[29\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08741_ _08749_/CLK line[67] VGND VGND VPWR VPWR _08741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05953_ _05929_/CLK line[73] VGND VGND VPWR VPWR _05953_/Q sky130_fd_sc_hd__dfxtp_1
X_08672_ _08672_/A _08687_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_05884_ _05884_/A _05887_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05752__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07623_ _07633_/CLK line[68] VGND VGND VPWR VPWR _07623_/Q sky130_fd_sc_hd__dfxtp_1
X_07554_ _07553_/Q _07567_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12585__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06505_ _06489_/CLK line[69] VGND VGND VPWR VPWR _06505_/Q sky130_fd_sc_hd__dfxtp_1
X_07485_ _07467_/CLK line[5] VGND VGND VPWR VPWR _07486_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[16\].CGAND _07111_/A wr VGND VGND VPWR VPWR OVHB\[16\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__07679__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09224_ _09223_/Q _09247_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06583__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07041__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06436_ _06435_/Q _06447_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06367_ _06353_/CLK line[6] VGND VGND VPWR VPWR _06368_/A sky130_fd_sc_hd__dfxtp_1
X_09155_ _09147_/CLK line[15] VGND VGND VPWR VPWR _09155_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].CG clk OVHB\[0\].CG/GATE VGND VGND VPWR VPWR OVHB\[0\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_120_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09894__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08106_ _08105_/Q _08127_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_05318_ _05317_/Q _05327_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_06298_ _06297_/Q _06307_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_09086_ _09086_/A _09107_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VALID\[12\].FF OVHB\[19\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[19\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05249_ _05253_/CLK line[7] VGND VGND VPWR VPWR _05249_/Q sky130_fd_sc_hd__dfxtp_1
X_08037_ _08033_/CLK line[1] VGND VGND VPWR VPWR _08037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10833__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05927__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08303__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09988_ _09987_/Q _10017_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08939_ _08947_/CLK line[44] VGND VGND VPWR VPWR _08940_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06758__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07216__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ _11949_/Q _11977_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09134__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10901_ _10903_/CLK line[45] VGND VGND VPWR VPWR _10902_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[22\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _11901_/CLK line[109] VGND VGND VPWR VPWR _11881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[15\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13620_ _13620_/CLK _13621_/X VGND VGND VPWR VPWR _13598_/CLK sky130_fd_sc_hd__dlclkp_1
X_10832_ _10832_/A _10857_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_13551_ _13552_/A wr VGND VGND VPWR VPWR _13551_/X sky130_fd_sc_hd__and2_1
X_10763_ _10783_/CLK line[110] VGND VGND VPWR VPWR _10763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].CGAND_A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DECH.DEC0.AND3_B A_h[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12502_ _13943_/X VGND VGND VPWR VPWR _12502_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06493__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13482_ _13552_/A VGND VGND VPWR VPWR _13482_/Y sky130_fd_sc_hd__inv_2
X_10694_ _10693_/Q _10717_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12433_ _12449_/CLK line[96] VGND VGND VPWR VPWR _12433_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[11\].TOBUF OVHB\[19\].VALID\[11\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12364_ _12363_/Q _12397_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_11315_ _11343_/CLK line[106] VGND VGND VPWR VPWR _11315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12295_ _12311_/CLK line[42] VGND VGND VPWR VPWR _12295_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09309__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11246_ _11246_/A _11277_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11177_ _11191_/CLK line[43] VGND VGND VPWR VPWR _11178_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10128_ _10127_/Q _10157_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11574__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10059_ _10073_/CLK line[44] VGND VGND VPWR VPWR _10059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06668__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09044__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11871__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[20\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08883__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13818_ _13822_/CLK line[84] VGND VGND VPWR VPWR _13818_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[10\].TOBUF OVHB\[12\].VALID\[10\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_13749_ _13748_/Q _13762_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07270_ _07269_/Q _07287_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].VALID\[10\].FF OVHB\[1\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[1\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06221_ _06223_/CLK line[67] VGND VGND VPWR VPWR _06221_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06152_ _06151_/Q _06167_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[19\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _07880_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11749__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05103_ _05093_/CLK line[68] VGND VGND VPWR VPWR _05103_/Q sky130_fd_sc_hd__dfxtp_1
X_06083_ _06077_/CLK line[4] VGND VGND VPWR VPWR _06083_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09219__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05034_ _05033_/Q _05047_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_09911_ _09912_/A wr VGND VGND VPWR VPWR _09911_/X sky130_fd_sc_hd__and2_1
XANTENNA__08123__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09842_ _09912_/A VGND VGND VPWR VPWR _09842_/Y sky130_fd_sc_hd__inv_2
X_09773_ _09793_/CLK line[32] VGND VGND VPWR VPWR _09773_/Q sky130_fd_sc_hd__dfxtp_1
X_06985_ _07001_/CLK line[47] VGND VGND VPWR VPWR _06986_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[1\].FF OVHB\[8\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[8\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08724_ _08723_/Q _08757_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05936_ _05935_/Q _05957_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05482__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08655_ _08663_/CLK line[42] VGND VGND VPWR VPWR _08655_/Q sky130_fd_sc_hd__dfxtp_1
X_05867_ _05871_/CLK line[33] VGND VGND VPWR VPWR _05868_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08793__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07606_ _07605_/Q _07637_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08586_ _08585_/Q _08617_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_05798_ _05797_/Q _05817_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _07539_/CLK line[43] VGND VGND VPWR VPWR _07537_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07987__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07468_ _07467_/Q _07497_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09207_ _09206_/Q _09212_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_06419_ _06421_/CLK line[44] VGND VGND VPWR VPWR _06419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07399_ _07393_/CLK line[108] VGND VGND VPWR VPWR _07399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09138_ _09116_/CLK line[121] VGND VGND VPWR VPWR _09138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10563__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09069_ _09069_/A _09072_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05657__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11100_ _11100_/CLK _11101_/X VGND VGND VPWR VPWR _11090_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.MUX\[0\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08033__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12080_ _12080_/CLK _12081_/X VGND VGND VPWR VPWR _12072_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13874__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11031_ _11032_/A wr VGND VGND VPWR VPWR _11031_/X sky130_fd_sc_hd__and2_1
XANTENNA__08968__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[18\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _07495_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07872__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06131__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[9\].VALID\[9\].TOBUF OVHB\[9\].VALID\[9\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ _12962_/CLK line[86] VGND VGND VPWR VPWR _12982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11933_ _11933_/A _11942_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09799__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11864_ _11846_/CLK line[87] VGND VGND VPWR VPWR _11864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[30\].CGAND_A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13603_ _13602_/Q _13622_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_10815_ _10814_/Q _10822_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10738__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[10\].FF OVHB\[15\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[15\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[3\].FF OVHB\[6\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[6\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11795_ _11795_/A _11802_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13114__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13534_ _13528_/CLK line[82] VGND VGND VPWR VPWR _13535_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08208__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10746_ _10728_/CLK line[88] VGND VGND VPWR VPWR _10746_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12953__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13411__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13465_ _13464_/Q _13482_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_10677_ _10676_/Q _10682_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_12416_ _12414_/CLK line[83] VGND VGND VPWR VPWR _12416_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06306__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13396_ _13394_/CLK line[19] VGND VGND VPWR VPWR _13396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10473__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12347_ _12346_/Q _12362_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[4\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12278_ _12268_/CLK line[20] VGND VGND VPWR VPWR _12279_/A sky130_fd_sc_hd__dfxtp_1
X_11229_ _11229_/A _11242_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07782__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06398__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06770_ _06770_/A _06797_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09352__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05721_ _05739_/CLK line[109] VGND VGND VPWR VPWR _05721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08440_ _08440_/CLK _08441_/X VGND VGND VPWR VPWR _08410_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09071__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05652_ _05651_/Q _05677_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10648__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05583_ _05575_/CLK line[46] VGND VGND VPWR VPWR _05583_/Q sky130_fd_sc_hd__dfxtp_1
X_08371_ _13921_/X wr VGND VGND VPWR VPWR _08371_/X sky130_fd_sc_hd__and2_1
XOVHB\[16\].VALID\[4\].TOBUF OVHB\[16\].VALID\[4\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_07322_ _13918_/X VGND VGND VPWR VPWR _07322_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07022__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07253_ _07267_/CLK line[32] VGND VGND VPWR VPWR _07253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12863__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07957__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06861__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06204_ _06203_/Q _06237_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_07184_ _07183_/Q _07217_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11479__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[5\].FF OVHB\[4\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[4\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06135_ _06147_/CLK line[42] VGND VGND VPWR VPWR _06136_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10961__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09527__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06066_ _06065_/Q _06097_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05017_ _05041_/CLK line[43] VGND VGND VPWR VPWR _05017_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[23\]_A2 _06545_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09246__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08788__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09825_ _09825_/A _09842_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12103__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09756_ _09760_/CLK line[19] VGND VGND VPWR VPWR _09756_/Q sky130_fd_sc_hd__dfxtp_1
X_06968_ _06960_/CLK line[25] VGND VGND VPWR VPWR _06969_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08707_ _08707_/A _08722_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05919_ _05918_/Q _05922_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09687_ _09686_/Q _09702_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_06899_ _06898_/Q _06902_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_08638_ _08646_/CLK line[20] VGND VGND VPWR VPWR _08638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09412__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08569_ _08569_/A _08582_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _10594_/CLK line[21] VGND VGND VPWR VPWR _10600_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _11588_/CLK line[85] VGND VGND VPWR VPWR _11580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10531_ _10530_/Q _10542_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06771__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13250_ _13254_/CLK line[95] VGND VGND VPWR VPWR _13250_/Q sky130_fd_sc_hd__dfxtp_1
X_10462_ _10466_/CLK line[86] VGND VGND VPWR VPWR _10462_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11389__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12201_ _12200_/Q _12222_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10293__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13181_ _13181_/A _13202_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_10393_ _10393_/A _10402_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05387__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12132_ _12130_/CLK line[81] VGND VGND VPWR VPWR _12133_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[3\].TOBUF OVHB\[22\].VALID\[3\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__08698__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12063_ _12062_/Q _12082_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_11014_ _11002_/CLK line[82] VGND VGND VPWR VPWR _11014_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[7\].FF OVHB\[2\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[2\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12013__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06796__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06011__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12965_ _12964_/Q _12992_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11852__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11207__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11916_ _11934_/CLK line[125] VGND VGND VPWR VPWR _11916_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06946__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12896_ _12902_/CLK line[61] VGND VGND VPWR VPWR _12896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09322__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10468__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11847_ _11847_/A _11872_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[17\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XMUX.MUX\[2\] _09160_/Z _05030_/Z _06780_/Z _13570_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[2] sky130_fd_sc_hd__mux4_1
X_11778_ _11776_/CLK line[62] VGND VGND VPWR VPWR _11778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13779__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13517_ _13552_/A VGND VGND VPWR VPWR _13517_/Y sky130_fd_sc_hd__inv_2
X_10729_ _10728_/Q _10752_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_13448_ _13468_/CLK line[48] VGND VGND VPWR VPWR _13448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13379_ _13378_/Q _13412_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05297__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07940_ _07946_/CLK line[85] VGND VGND VPWR VPWR _07941_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[1\].FF OVHB\[30\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[30\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[31\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08401__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[9\].TOBUF OVHB\[14\].VALID\[9\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_07871_ _07870_/Q _07882_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13019__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09610_ _09626_/CLK line[95] VGND VGND VPWR VPWR _09610_/Q sky130_fd_sc_hd__dfxtp_1
X_06822_ _06802_/CLK line[86] VGND VGND VPWR VPWR _06822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12501__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09541_ _09540_/Q _09562_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_06753_ _06752_/Q _06762_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05704_ _05708_/CLK line[87] VGND VGND VPWR VPWR _05704_/Q sky130_fd_sc_hd__dfxtp_1
X_09472_ _09482_/CLK line[17] VGND VGND VPWR VPWR _09473_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05760__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06684_ _06682_/CLK line[23] VGND VGND VPWR VPWR _06685_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[9\].FF OVHB\[0\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[0\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ _08422_/Q _08442_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10378__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05635_ _05635_/A _05642_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _08358_/CLK line[18] VGND VGND VPWR VPWR _08355_/A sky130_fd_sc_hd__dfxtp_1
X_05566_ _05568_/CLK line[24] VGND VGND VPWR VPWR _05567_/A sky130_fd_sc_hd__dfxtp_1
X_07305_ _07305_/A _07322_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12593__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05497_ _05497_/A _05502_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_08285_ _08284_/Q _08302_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[13\].TOBUF OVHB\[9\].VALID\[13\].FF/Q OVHB\[9\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07687__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07236_ _07232_/CLK line[19] VGND VGND VPWR VPWR _07236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07167_ _07166_/Q _07182_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11002__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06118_ _06108_/CLK line[20] VGND VGND VPWR VPWR _06118_/Q sky130_fd_sc_hd__dfxtp_1
X_07098_ _07098_/CLK line[84] VGND VGND VPWR VPWR _07099_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[2\].FF OVHB\[29\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[29\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08161__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05000__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10841__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06049_ _06048_/Q _06062_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05935__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08311__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09808_ _09834_/CLK line[48] VGND VGND VPWR VPWR _09809_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12768__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09739_ _09738_/Q _09772_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04934__B1 A_h[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12750_ _12774_/CLK line[122] VGND VGND VPWR VPWR _12750_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[12\].TOBUF OVHB\[2\].VALID\[12\].FF/Q OVHB\[2\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11700_/Q _11732_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12681_ _12681_/A _12712_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[8\].TOBUF OVHB\[20\].VALID\[8\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11636_/CLK line[123] VGND VGND VPWR VPWR _11632_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08336__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _11562_/Q _11592_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ _13301_/Q _13307_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ _10520_/CLK line[124] VGND VGND VPWR VPWR _10514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ _11500_/CLK line[60] VGND VGND VPWR VPWR _11494_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11697__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13233_ _13213_/CLK line[73] VGND VGND VPWR VPWR _13233_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12008__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10445_ _10445_/A _10472_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13164_ _13164_/A _13167_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10376_ _10384_/CLK line[61] VGND VGND VPWR VPWR _10376_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _13795_/CLK sky130_fd_sc_hd__clkbuf_4
X_12115_ _12115_/CLK _12116_/X VGND VGND VPWR VPWR _12109_/CLK sky130_fd_sc_hd__dlclkp_1
X_13095_ _13095_/CLK _13096_/X VGND VGND VPWR VPWR _13075_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_2_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12046_ _12151_/A wr VGND VGND VPWR VPWR _12046_/X sky130_fd_sc_hd__and2_1
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[27\].VALID\[4\].FF OVHB\[27\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[27\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12678__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11582__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[5\]_A2 _13506_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06676__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[10\].FF OVHB\[6\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[6\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12948_ _12947_/Q _12957_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09052__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12879_ _12881_/CLK line[39] VGND VGND VPWR VPWR _12879_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09987__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08891__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05420_ _05424_/CLK line[85] VGND VGND VPWR VPWR _05420_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[13\]_A1 _05582_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05351_ _05350_/Q _05362_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12991__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05282_ _05278_/CLK line[22] VGND VGND VPWR VPWR _05282_/Q sky130_fd_sc_hd__dfxtp_1
X_08070_ _08070_/CLK line[31] VGND VGND VPWR VPWR _08070_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07300__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07021_ _07020_/Q _07042_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[15\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11757__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[4\].VALID\[0\].TOBUF OVHB\[4\].VALID\[0\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08972_ _08972_/CLK line[59] VGND VGND VPWR VPWR _08972_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10016__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09227__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07923_ _07922_/Q _07952_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[3\].TOBUF OVHB\[29\].VALID\[3\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XDATA\[8\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _13410_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_99_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07854_ _07854_/CLK line[60] VGND VGND VPWR VPWR _07855_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06805_ _06804_/Q _06832_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04916__B1 _04916_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11492__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07785_ _07784_/Q _07812_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_04997_ _04996_/Q _05012_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_09524_ _09523_/Q _09527_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_06736_ _06740_/CLK line[61] VGND VGND VPWR VPWR _06736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05490__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[8\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09455_ _09455_/CLK _09456_/X VGND VGND VPWR VPWR _09427_/CLK sky130_fd_sc_hd__dlclkp_1
X_06667_ _06667_/A _06692_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ _13921_/X wr VGND VGND VPWR VPWR _08406_/X sky130_fd_sc_hd__and2_1
XANTENNA__13062__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05618_ _05632_/CLK line[62] VGND VGND VPWR VPWR _05618_/Q sky130_fd_sc_hd__dfxtp_1
X_09386_ _09352_/A wr VGND VGND VPWR VPWR _09386_/X sky130_fd_sc_hd__and2_1
XFILLER_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[25\].VALID\[6\].FF OVHB\[25\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[25\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[14\].TOBUF OVHB\[25\].VALID\[14\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_06598_ _06596_/CLK line[126] VGND VGND VPWR VPWR _06599_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08337_ _13921_/X VGND VGND VPWR VPWR _08337_/Y sky130_fd_sc_hd__inv_2
X_05549_ _05548_/Q _05572_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08268_ _08282_/CLK line[112] VGND VGND VPWR VPWR _08268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07219_ _07218_/Q _07252_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_08199_ _08198_/Q _08232_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _10248_/CLK line[122] VGND VGND VPWR VPWR _10230_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[28\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _10750_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11667__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10571__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10161_ _10160_/Q _10192_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05665__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08041__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10092_ _10100_/CLK line[59] VGND VGND VPWR VPWR _10092_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13882__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13237__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08976__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13920_ _13923_/C _13923_/B _13922_/B _13923_/D VGND VGND VPWR VPWR _13920_/X sky130_fd_sc_hd__and4b_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13851_ _13845_/CLK line[99] VGND VGND VPWR VPWR _13852_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12498__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _12801_/Q _12817_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13782_ _13781_/Q _13797_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10994_ _10993_/Q _10997_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_12733_ _12741_/CLK line[100] VGND VGND VPWR VPWR _12734_/A sky130_fd_sc_hd__dfxtp_1
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12664_/A _12677_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09600__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11605_/CLK line[101] VGND VGND VPWR VPWR _11615_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10746__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12601_/CLK line[37] VGND VGND VPWR VPWR _12596_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13122__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _11545_/Q _11557_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08216__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11477_ _11479_/CLK line[38] VGND VGND VPWR VPWR _11477_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[8\].FF OVHB\[23\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[23\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13216_ _13215_/Q _13237_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_10428_ _10427_/Q _10437_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10481__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13147_ _13163_/CLK line[33] VGND VGND VPWR VPWR _13147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10359_ _10341_/CLK line[39] VGND VGND VPWR VPWR _10360_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05575__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13078_ _13078_/A _13097_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[27\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _10365_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04920_ A_h[22] _04920_/B2 A_h[22] _04920_/B2 VGND VGND VPWR VPWR _04921_/D sky130_fd_sc_hd__a2bb2o_4
X_12029_ _12019_/CLK line[34] VGND VGND VPWR VPWR _12029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07790__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[31\].INV _13979_/X VGND VGND VPWR VPWR OVHB\[31\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_81_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07570_ _07572_/CLK line[58] VGND VGND VPWR VPWR _07570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06521_ _06520_/Q _06552_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _09240_/A _09247_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_06452_ _06464_/CLK line[59] VGND VGND VPWR VPWR _06453_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[5\].TOBUF OVHB\[2\].VALID\[5\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_05403_ _05402_/Q _05432_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10656__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09171_ _09147_/CLK line[8] VGND VGND VPWR VPWR _09171_/Q sky130_fd_sc_hd__dfxtp_1
X_06383_ _06382_/Q _06412_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13032__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[8\].TOBUF OVHB\[27\].VALID\[8\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_08122_ _08121_/Q _08127_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_05334_ _05332_/CLK line[60] VGND VGND VPWR VPWR _05334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07030__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12871__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08053_ _08033_/CLK line[9] VGND VGND VPWR VPWR _08053_/Q sky130_fd_sc_hd__dfxtp_1
X_05265_ _05264_/Q _05292_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07965__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07004_ _07004_/A _07007_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_05196_ _05214_/CLK line[125] VGND VGND VPWR VPWR _05196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[12\].CGAND _13910_/X wr VGND VGND VPWR VPWR OVHB\[12\].CGAND/X sky130_fd_sc_hd__and2_4
X_08955_ _08947_/CLK line[37] VGND VGND VPWR VPWR _08955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[13\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07906_ _07905_/Q _07917_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08886_ _08885_/Q _08897_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07837_ _07837_/CLK line[38] VGND VGND VPWR VPWR _07838_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13207__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12111__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07768_ _07767_/Q _07777_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07205__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09507_ _09507_/CLK line[33] VGND VGND VPWR VPWR _09508_/A sky130_fd_sc_hd__dfxtp_1
X_06719_ _06711_/CLK line[39] VGND VGND VPWR VPWR _06719_/Q sky130_fd_sc_hd__dfxtp_1
X_07699_ _07679_/CLK line[103] VGND VGND VPWR VPWR _07700_/A sky130_fd_sc_hd__dfxtp_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[16\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _07110_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09457_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XMUX.MUX\[20\] _10039_/Z _13469_/Z _06539_/Z _07169_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[20] sky130_fd_sc_hd__mux4_1
XFILLER_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09369_ _09365_/CLK line[98] VGND VGND VPWR VPWR _09370_/A sky130_fd_sc_hd__dfxtp_1
X_11400_ _11400_/A _11417_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12380_ _12379_/Q _12397_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11331_ _11343_/CLK line[99] VGND VGND VPWR VPWR _11332_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11262_ _11261_/Q _11277_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11397__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13001_ _12999_/CLK line[109] VGND VGND VPWR VPWR _13001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10213_ _10217_/CLK line[100] VGND VGND VPWR VPWR _10213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11193_ _11191_/CLK line[36] VGND VGND VPWR VPWR _11193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10144_ _10143_/Q _10157_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10075_ _10073_/CLK line[37] VGND VGND VPWR VPWR _10075_/Q sky130_fd_sc_hd__dfxtp_1
X_13903_ A[4] VGND VGND VPWR VPWR _13909_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12021__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13834_ _13833_/Q _13867_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07115__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[30\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ _13763_/CLK line[74] VGND VGND VPWR VPWR _13765_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11860__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10977_ _10977_/CLK line[65] VGND VGND VPWR VPWR _10978_/A sky130_fd_sc_hd__dfxtp_1
X_12716_ _12715_/Q _12747_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06954__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13696_ _13695_/Q _13727_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09330__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ _12667_/CLK line[75] VGND VGND VPWR VPWR _12647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[23\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[15\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _06725_/CLK sky130_fd_sc_hd__clkbuf_4
X_12578_ _12577_/Q _12607_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13787__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11529_ _11535_/CLK line[76] VGND VGND VPWR VPWR _11530_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12046__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05050_ _05058_/CLK line[58] VGND VGND VPWR VPWR _05050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[16\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08740_ _08739_/Q _08757_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_05952_ _05952_/A _05957_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09505__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08671_ _08663_/CLK line[35] VGND VGND VPWR VPWR _08672_/A sky130_fd_sc_hd__dfxtp_1
X_05883_ _05871_/CLK line[41] VGND VGND VPWR VPWR _05884_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07622_ _07621_/Q _07637_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_07553_ _07539_/CLK line[36] VGND VGND VPWR VPWR _07553_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06504_ _06503_/Q _06517_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07484_ _07483_/Q _07497_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_09223_ _09241_/CLK line[46] VGND VGND VPWR VPWR _09223_/Q sky130_fd_sc_hd__dfxtp_1
X_06435_ _06421_/CLK line[37] VGND VGND VPWR VPWR _06435_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10386__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09154_ _09153_/Q _09177_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_06366_ _06365_/Q _06377_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13697__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08105_ _08113_/CLK line[47] VGND VGND VPWR VPWR _08105_/Q sky130_fd_sc_hd__dfxtp_1
X_05317_ _05299_/CLK line[38] VGND VGND VPWR VPWR _05317_/Q sky130_fd_sc_hd__dfxtp_1
X_09085_ _09085_/CLK line[111] VGND VGND VPWR VPWR _09086_/A sky130_fd_sc_hd__dfxtp_1
X_06297_ _06285_/CLK line[102] VGND VGND VPWR VPWR _06297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07695__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VOBUF OVHB\[6\].V/Q OVHB\[6\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_08036_ _08035_/Q _08057_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_05248_ _05247_/Q _05257_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[26\]_A0 _11421_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[27\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11010__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05179_ _05157_/CLK line[103] VGND VGND VPWR VPWR _05179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06104__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09987_ _10011_/CLK line[11] VGND VGND VPWR VPWR _09987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11945__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08938_ _08937_/Q _08967_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05943__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08869_ _08869_/CLK line[12] VGND VGND VPWR VPWR _08869_/Q sky130_fd_sc_hd__dfxtp_1
X_10900_ _10899_/Q _10927_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_11880_ _11880_/A _11907_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10831_ _10843_/CLK line[13] VGND VGND VPWR VPWR _10832_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12776__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[15\].VALID\[12\].TOBUF OVHB\[15\].VALID\[12\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_13550_ _13550_/CLK _13551_/X VGND VGND VPWR VPWR _13528_/CLK sky130_fd_sc_hd__dlclkp_1
X_10762_ _10761_/Q _10787_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_12501_ _13943_/X wr VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[19\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13481_ _13552_/A wr VGND VGND VPWR VPWR _13481_/X sky130_fd_sc_hd__and2_1
XFILLER_13_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10693_ _10707_/CLK line[78] VGND VGND VPWR VPWR _10693_/Q sky130_fd_sc_hd__dfxtp_1
X_12432_ _13943_/X VGND VGND VPWR VPWR _12432_/Y sky130_fd_sc_hd__inv_2
XOVHB\[9\].VALID\[5\].TOBUF OVHB\[9\].VALID\[5\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12363_ _12387_/CLK line[64] VGND VGND VPWR VPWR _12363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13400__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11314_ _11313_/Q _11347_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12294_ _12293_/Q _12327_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[1\].INV _13984_/X VGND VGND VPWR VPWR OVHB\[1\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_49_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11245_ _11251_/CLK line[74] VGND VGND VPWR VPWR _11246_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ _11175_/Q _11207_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10127_ _10145_/CLK line[75] VGND VGND VPWR VPWR _10127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[0\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05853__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10058_ _10057_/Q _10087_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13817_ _13816_/Q _13832_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12686__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06684__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ _13746_/CLK line[52] VGND VGND VPWR VPWR _13748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09060__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13679_ _13678_/Q _13692_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09995__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06220_ _06219_/Q _06237_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_06151_ _06147_/CLK line[35] VGND VGND VPWR VPWR _06151_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10934__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13310__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05102_ _05101_/Q _05117_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_06082_ _06081_/Q _06097_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_05033_ _05041_/CLK line[36] VGND VGND VPWR VPWR _05033_/Q sky130_fd_sc_hd__dfxtp_1
X_09910_ _09910_/CLK _09911_/X VGND VGND VPWR VPWR _09908_/CLK sky130_fd_sc_hd__dlclkp_1
X_09841_ _09912_/A wr VGND VGND VPWR VPWR _09841_/X sky130_fd_sc_hd__and2_1
XOVHB\[16\].VALID\[0\].TOBUF OVHB\[16\].VALID\[0\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06859__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09772_ _09912_/A VGND VGND VPWR VPWR _09772_/Y sky130_fd_sc_hd__inv_2
X_06984_ _06983_/Q _07007_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09235__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08723_ _08749_/CLK line[64] VGND VGND VPWR VPWR _08723_/Q sky130_fd_sc_hd__dfxtp_1
X_05935_ _05929_/CLK line[79] VGND VGND VPWR VPWR _05935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08654_ _08653_/Q _08687_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_05866_ _05865_/Q _05887_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_07605_ _07633_/CLK line[74] VGND VGND VPWR VPWR _07605_/Q sky130_fd_sc_hd__dfxtp_1
X_08585_ _08609_/CLK line[10] VGND VGND VPWR VPWR _08585_/Q sky130_fd_sc_hd__dfxtp_1
X_05797_ _05799_/CLK line[1] VGND VGND VPWR VPWR _05797_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07536_ _07535_/Q _07567_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06594__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07467_ _07467_/CLK line[11] VGND VGND VPWR VPWR _07467_/Q sky130_fd_sc_hd__dfxtp_1
X_09206_ _09200_/CLK line[24] VGND VGND VPWR VPWR _09206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06418_ _06417_/Q _06447_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_07398_ _07397_/Q _07427_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09137_ _09136_/Q _09142_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_06349_ _06353_/CLK line[12] VGND VGND VPWR VPWR _06349_/Q sky130_fd_sc_hd__dfxtp_1
X_09068_ _09068_/CLK line[89] VGND VGND VPWR VPWR _09069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08019_ _08018_/Q _08022_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[0\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11030_ _11030_/CLK _11031_/X VGND VGND VPWR VPWR _11002_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06412__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11675__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06769__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05673__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06131__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09145__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12981_ _12980_/Q _12992_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13890__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08984__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _11934_/CLK line[118] VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11863_ _11862_/Q _11872_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10814_ _10804_/CLK line[119] VGND VGND VPWR VPWR _10814_/Q sky130_fd_sc_hd__dfxtp_1
X_13602_ _13598_/CLK line[113] VGND VGND VPWR VPWR _13602_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[30\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11794_ _11776_/CLK line[55] VGND VGND VPWR VPWR _11795_/A sky130_fd_sc_hd__dfxtp_1
X_13533_ _13533_/A _13552_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10745_ _10744_/Q _10752_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06009__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13464_ _13468_/CLK line[50] VGND VGND VPWR VPWR _13464_/Q sky130_fd_sc_hd__dfxtp_1
X_10676_ _10656_/CLK line[56] VGND VGND VPWR VPWR _10676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12415_ _12415_/A _12432_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_13395_ _13394_/Q _13412_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[8\].FF OVHB\[9\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[9\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06306__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05848__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12346_ _12352_/CLK line[51] VGND VGND VPWR VPWR _12346_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08224__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12277_ _12276_/Q _12292_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11228_ _11216_/CLK line[52] VGND VGND VPWR VPWR _11229_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11159_ _11158_/Q _11172_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05583__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[8\]_A0 _09452_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05720_ _05719_/Q _05747_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_05651_ _05671_/CLK line[77] VGND VGND VPWR VPWR _05651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08370_ _08370_/CLK _08371_/X VGND VGND VPWR VPWR _08358_/CLK sky130_fd_sc_hd__dlclkp_1
X_05582_ _05581_/Q _05607_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07321_ _13918_/X wr VGND VGND VPWR VPWR _07321_/X sky130_fd_sc_hd__and2_1
XDATA\[6\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _13025_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[14\].VALID\[5\].TOBUF OVHB\[14\].VALID\[5\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07252_ _13918_/X VGND VGND VPWR VPWR _07252_/Y sky130_fd_sc_hd__inv_2
X_06203_ _06223_/CLK line[64] VGND VGND VPWR VPWR _06203_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10664__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07183_ _07183_/CLK line[0] VGND VGND VPWR VPWR _07183_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13040__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05758__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06134_ _06133_/Q _06167_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08134__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10961__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06065_ _06077_/CLK line[10] VGND VGND VPWR VPWR _06065_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[31\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07973__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05016_ _05015_/Q _05047_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_MUX.MUX\[23\]_A3 _09415_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09824_ _09834_/CLK line[50] VGND VGND VPWR VPWR _09825_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06967_ _06966_/Q _06972_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_09755_ _09754_/Q _09772_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08706_ _08710_/CLK line[51] VGND VGND VPWR VPWR _08707_/A sky130_fd_sc_hd__dfxtp_1
X_05918_ _05902_/CLK line[57] VGND VGND VPWR VPWR _05918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09686_ _09694_/CLK line[115] VGND VGND VPWR VPWR _09686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06898_ _06892_/CLK line[121] VGND VGND VPWR VPWR _06898_/Q sky130_fd_sc_hd__dfxtp_1
X_08637_ _08636_/Q _08652_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10839__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05849_ _05848_/Q _05852_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13215__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08568_ _08560_/CLK line[116] VGND VGND VPWR VPWR _08569_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07213__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07519_ _07518_/Q _07532_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _08498_/Q _08512_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _10520_/CLK line[117] VGND VGND VPWR VPWR _10530_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A _10472_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[5\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _12640_/CLK sky130_fd_sc_hd__clkbuf_4
X_12200_ _12204_/CLK line[127] VGND VGND VPWR VPWR _12200_/Q sky130_fd_sc_hd__dfxtp_1
X_13180_ _13194_/CLK line[63] VGND VGND VPWR VPWR _13181_/A sky130_fd_sc_hd__dfxtp_1
X_10392_ _10384_/CLK line[54] VGND VGND VPWR VPWR _10393_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[0\].FF OVHB\[18\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[18\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12131_ _12131_/A _12152_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07883__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12062_ _12072_/CLK line[49] VGND VGND VPWR VPWR _12062_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[4\].TOBUF OVHB\[20\].VALID\[4\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_11013_ _11012_/Q _11032_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06499__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06796__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12964_ _12962_/CLK line[92] VGND VGND VPWR VPWR _12964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11915_ _11914_/Q _11942_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_12895_ _12894_/Q _12922_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11846_ _11846_/CLK line[93] VGND VGND VPWR VPWR _11847_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07123__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12964__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[25\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _09980_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[23\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _11776_/Q _11802_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_13516_ _13552_/A wr VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__and2_1
X_10728_ _10728_/CLK line[94] VGND VGND VPWR VPWR _10728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06962__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05221__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10659_ _10659_/A _10682_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
X_13447_ _13552_/A VGND VGND VPWR VPWR _13447_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13378_ _13394_/CLK line[16] VGND VGND VPWR VPWR _13378_/Q sky130_fd_sc_hd__dfxtp_1
X_12329_ _12328_/Q _12362_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08889__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[4\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _12255_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07870_ _07854_/CLK line[53] VGND VGND VPWR VPWR _07870_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12204__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[2\].FF OVHB\[16\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[16\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06821_ _06820_/Q _06832_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12501__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09540_ _09554_/CLK line[63] VGND VGND VPWR VPWR _09540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06752_ _06740_/CLK line[54] VGND VGND VPWR VPWR _06752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09513__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05703_ _05703_/A _05712_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09471_ _09470_/Q _09492_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[14\].TOBUF OVHB\[5\].VALID\[14\].FF/Q OVHB\[5\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_58_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06683_ _06682_/Q _06692_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_08422_ _08410_/CLK line[49] VGND VGND VPWR VPWR _08422_/Q sky130_fd_sc_hd__dfxtp_1
X_05634_ _05632_/CLK line[55] VGND VGND VPWR VPWR _05635_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[17\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08353_ _08352_/Q _08372_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].V OVHB\[9\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[9\].V/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05565_ _05564_/Q _05572_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_07304_ _07292_/CLK line[50] VGND VGND VPWR VPWR _07305_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06872__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08284_ _08282_/CLK line[114] VGND VGND VPWR VPWR _08284_/Q sky130_fd_sc_hd__dfxtp_1
X_05496_ _05476_/CLK line[120] VGND VGND VPWR VPWR _05497_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10394__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07235_ _07235_/A _07252_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05488__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[24\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _09595_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07166_ _07170_/CLK line[115] VGND VGND VPWR VPWR _07166_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08442__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06117_ _06116_/Q _06132_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08799__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04920__A1_N A_h[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07097_ _07096_/Q _07112_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08161__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06048_ _06050_/CLK line[116] VGND VGND VPWR VPWR _06048_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[10\].TOBUF OVHB\[25\].VALID\[10\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__04935__A1_N A_h[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09807_ _09912_/A VGND VGND VPWR VPWR _09807_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06112__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07999_ _07998_/Q _08022_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11953__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09738_ _09760_/CLK line[16] VGND VGND VPWR VPWR _09738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04934__B2 _04934_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05951__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09423__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10569__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09668_/Q _09702_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11706_/CLK line[26] VGND VGND VPWR VPWR _11700_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08039__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12680_ _12708_/CLK line[90] VGND VGND VPWR VPWR _12681_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[14\].VALID\[4\].FF OVHB\[14\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[14\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11631_ _11630_/Q _11662_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[8\].FF OVHB\[31\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[31\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07878__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08336__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _11588_/CLK line[91] VGND VGND VPWR VPWR _11562_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13301_ _13285_/CLK line[104] VGND VGND VPWR VPWR _13301_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _10512_/Q _10542_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _11492_/Q _11522_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05398__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13232_ _13231_/Q _13237_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_10444_ _10466_/CLK line[92] VGND VGND VPWR VPWR _10445_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13163_ _13163_/CLK line[41] VGND VGND VPWR VPWR _13164_/A sky130_fd_sc_hd__dfxtp_1
X_10375_ _10374_/Q _10402_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _12113_/Q _12117_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08502__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[23\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _09210_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_2_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13094_ _13093_/Q _13097_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12045_ _12045_/CLK _12046_/X VGND VGND VPWR VPWR _12019_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[23\].V OVHB\[23\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[23\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[13\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _06340_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_120_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04925__A1 A_h[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10122__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04925__B2 _04923_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05861__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09911__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10479__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[5\]_A3 _05176_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12947_ _12937_/CLK line[70] VGND VGND VPWR VPWR _12947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12878_ _12877_/Q _12887_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12694__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11829_ _11823_/CLK line[71] VGND VGND VPWR VPWR _11829_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[13\]_A2 _10972_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07788__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05350_ _05332_/CLK line[53] VGND VGND VPWR VPWR _05350_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12991__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05281_ _05280_/Q _05292_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11103__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07020_ _07030_/CLK line[63] VGND VGND VPWR VPWR _07020_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[6\].FF OVHB\[12\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[12\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05886__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[21\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05101__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10942__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08412__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08971_ _08970_/Q _09002_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10016__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[1\].TOBUF OVHB\[2\].VALID\[1\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_07922_ _07946_/CLK line[91] VGND VGND VPWR VPWR _07922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[14\].V OVHB\[14\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[14\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07028__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[4\].TOBUF OVHB\[27\].VALID\[4\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_07853_ _07852_/Q _07882_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12869__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06804_ _06802_/CLK line[92] VGND VGND VPWR VPWR _06804_/Q sky130_fd_sc_hd__dfxtp_1
X_07784_ _07788_/CLK line[28] VGND VGND VPWR VPWR _07784_/Q sky130_fd_sc_hd__dfxtp_1
X_04996_ _05000_/CLK line[19] VGND VGND VPWR VPWR _04996_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09243__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06735_ _06734_/Q _06762_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_09523_ _09507_/CLK line[41] VGND VGND VPWR VPWR _09523_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[12\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _05955_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_65_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09454_ _09453_/Q _09457_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_06666_ _06682_/CLK line[29] VGND VGND VPWR VPWR _06667_/A sky130_fd_sc_hd__dfxtp_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05617_ _05616_/Q _05642_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_08405_ _08405_/CLK _08406_/X VGND VGND VPWR VPWR _08383_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_52_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09385_ _09385_/CLK _09386_/X VGND VGND VPWR VPWR _09365_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_80_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06597_ _06597_/A _06622_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_08336_ _13921_/X wr VGND VGND VPWR VPWR _08336_/X sky130_fd_sc_hd__and2_1
X_05548_ _05568_/CLK line[30] VGND VGND VPWR VPWR _05548_/Q sky130_fd_sc_hd__dfxtp_1
X_08267_ _13940_/X VGND VGND VPWR VPWR _08267_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12109__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05479_ _05478_/Q _05502_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
X_07218_ _07232_/CLK line[16] VGND VGND VPWR VPWR _07218_/Q sky130_fd_sc_hd__dfxtp_1
X_08198_ _08208_/CLK line[80] VGND VGND VPWR VPWR _08198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07149_ _07148_/Q _07182_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09418__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _10188_/CLK line[90] VGND VGND VPWR VPWR _10160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10091_ _10090_/Q _10122_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[8\].FF OVHB\[10\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[10\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[11\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11683__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13850_ _13849_/Q _13867_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06777__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09153__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12801_ _12803_/CLK line[3] VGND VGND VPWR VPWR _12801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13781_ _13763_/CLK line[67] VGND VGND VPWR VPWR _13781_/Q sky130_fd_sc_hd__dfxtp_1
X_10993_ _10977_/CLK line[73] VGND VGND VPWR VPWR _10993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08992__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12732_ _12731_/Q _12747_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07251__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12667_/CLK line[68] VGND VGND VPWR VPWR _12664_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _05570_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11613_/Q _11627_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12594_/A _12607_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07401__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ _11535_/CLK line[69] VGND VGND VPWR VPWR _11545_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06017__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11476_ _11475_/Q _11487_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11858__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13215_ _13213_/CLK line[79] VGND VGND VPWR VPWR _13215_/Q sky130_fd_sc_hd__dfxtp_1
X_10427_ _10405_/CLK line[70] VGND VGND VPWR VPWR _10427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09328__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10358_ _10357_/Q _10367_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_13146_ _13145_/Q _13167_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13077_ _13075_/CLK line[1] VGND VGND VPWR VPWR _13078_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10289_ _10277_/CLK line[7] VGND VGND VPWR VPWR _10290_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12028_ _12027_/Q _12047_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07426__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11593__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05591__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13979_ _13979_/A _13979_/B _13979_/C _13979_/D VGND VGND VPWR VPWR _13979_/X sky130_fd_sc_hd__and4_4
XANTENNA__10787__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06520_ _06528_/CLK line[90] VGND VGND VPWR VPWR _06520_/Q sky130_fd_sc_hd__dfxtp_1
X_06451_ _06450_/Q _06482_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05402_ _05424_/CLK line[91] VGND VGND VPWR VPWR _05402_/Q sky130_fd_sc_hd__dfxtp_1
X_09170_ _09169_/Q _09177_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[6\].TOBUF OVHB\[0\].VALID\[6\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_06382_ _06408_/CLK line[27] VGND VGND VPWR VPWR _06382_/Q sky130_fd_sc_hd__dfxtp_1
X_08121_ _08113_/CLK line[40] VGND VGND VPWR VPWR _08121_/Q sky130_fd_sc_hd__dfxtp_1
X_05333_ _05332_/Q _05362_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[9\].TOBUF OVHB\[25\].VALID\[9\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_135_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08052_ _08052_/A _08057_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_05264_ _05278_/CLK line[28] VGND VGND VPWR VPWR _05264_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11768__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07003_ _07001_/CLK line[41] VGND VGND VPWR VPWR _07004_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10672__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05195_ _05194_/Q _05222_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05766__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08142__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[24\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08954_ _08953_/Q _08967_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07981__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12599__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07905_ _07905_/CLK line[69] VGND VGND VPWR VPWR _07905_/Q sky130_fd_sc_hd__dfxtp_1
X_08885_ _08869_/CLK line[5] VGND VGND VPWR VPWR _08885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07836_ _07835_/Q _07847_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VOBUF OVHB\[2\].V/Q OVHB\[2\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_07767_ _07773_/CLK line[6] VGND VGND VPWR VPWR _07767_/Q sky130_fd_sc_hd__dfxtp_1
X_04979_ _04978_/Q _05012_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11008__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09506_ _09505_/Q _09527_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06718_ _06718_/A _06727_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07698_ _07697_/Q _07707_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05006__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06649_ _06633_/CLK line[7] VGND VGND VPWR VPWR _06650_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10847__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09437_ _09427_/CLK line[1] VGND VGND VPWR VPWR _09438_/A sky130_fd_sc_hd__dfxtp_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13223__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08317__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09368_ _09367_/Q _09387_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[13\] _13352_/Z _05582_/Z _10972_/Z _13562_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[13] sky130_fd_sc_hd__mux4_1
XFILLER_36_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08319_ _08329_/CLK line[2] VGND VGND VPWR VPWR _08319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09299_ _09307_/CLK line[66] VGND VGND VPWR VPWR _09299_/Q sky130_fd_sc_hd__dfxtp_1
X_11330_ _11330_/A _11347_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[2\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10582__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _11251_/CLK line[67] VGND VGND VPWR VPWR _11261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10212_ _10212_/A _10227_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_13000_ _13000_/A _13027_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_11192_ _11191_/Q _11207_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10143_ _10145_/CLK line[68] VGND VGND VPWR VPWR _10143_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12152__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[8\].TOBUF OVHB\[31\].VALID\[8\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07891__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A _10087_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[1\].FF OVHB\[3\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[3\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[1\].TOBUF OVHB\[9\].VALID\[1\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_13902_ _13907_/X VGND VGND VPWR VPWR _13902_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13833_ _13845_/CLK line[96] VGND VGND VPWR VPWR _13833_/Q sky130_fd_sc_hd__dfxtp_1
X_13764_ _13763_/Q _13797_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A _10997_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_12715_ _12741_/CLK line[106] VGND VGND VPWR VPWR _12715_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10757__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13133__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13695_ _13701_/CLK line[42] VGND VGND VPWR VPWR _13695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _12645_/Q _12677_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12972__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12577_ _12601_/CLK line[43] VGND VGND VPWR VPWR _12577_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12327__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11527_/Q _11557_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12046__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11588__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11459_ _11479_/CLK line[44] VGND VGND VPWR VPWR _11460_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09058__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13129_ _13128_/Q _13132_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[25\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05951_ _05929_/CLK line[72] VGND VGND VPWR VPWR _05952_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13308__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[14\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08670_ _08670_/A _08687_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12212__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05882_ _05882_/A _05887_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07306__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07621_ _07633_/CLK line[67] VGND VGND VPWR VPWR _07621_/Q sky130_fd_sc_hd__dfxtp_1
X_07552_ _07552_/A _07567_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09521__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06503_ _06489_/CLK line[68] VGND VGND VPWR VPWR _06503_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[3\].FF OVHB\[1\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[1\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[14\].TOBUF OVHB\[18\].VALID\[14\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_07483_ _07467_/CLK line[4] VGND VGND VPWR VPWR _07483_/Q sky130_fd_sc_hd__dfxtp_1
X_09222_ _09222_/A _09247_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06434_ _06433_/Q _06447_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13621__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09153_ _09147_/CLK line[14] VGND VGND VPWR VPWR _09153_/Q sky130_fd_sc_hd__dfxtp_1
X_06365_ _06353_/CLK line[5] VGND VGND VPWR VPWR _06365_/Q sky130_fd_sc_hd__dfxtp_1
X_08104_ _08104_/A _08127_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_05316_ _05315_/Q _05327_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06880__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09084_ _09084_/A _09107_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06296_ _06296_/A _06307_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11498__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08035_ _08033_/CLK line[15] VGND VGND VPWR VPWR _08035_/Q sky130_fd_sc_hd__dfxtp_1
X_05247_ _05253_/CLK line[6] VGND VGND VPWR VPWR _05247_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05496__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[26\]_A1 _13451_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05178_ _05177_/Q _05187_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_09986_ _09985_/Q _10017_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08937_ _08947_/CLK line[43] VGND VGND VPWR VPWR _08937_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[13\].TOBUF OVHB\[11\].VALID\[13\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12122__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08868_ _08867_/Q _08897_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09281__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06120__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07819_ _07837_/CLK line[44] VGND VGND VPWR VPWR _07819_/Q sky130_fd_sc_hd__dfxtp_1
X_08799_ _08823_/CLK line[108] VGND VGND VPWR VPWR _08800_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11961__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].CGAND _13907_/X wr VGND VGND VPWR VPWR OVHB\[9\].CGAND/X sky130_fd_sc_hd__and2_4
X_10830_ _10829_/Q _10857_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09431__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ _10783_/CLK line[109] VGND VGND VPWR VPWR _10761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _12500_/CLK _12501_/X VGND VGND VPWR VPWR _12490_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08047__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13480_ _13480_/CLK _13481_/X VGND VGND VPWR VPWR _13468_/CLK sky130_fd_sc_hd__dlclkp_1
X_10692_ _10691_/Q _10717_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13888__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12431_ _13943_/X wr VGND VGND VPWR VPWR _12431_/X sky130_fd_sc_hd__and2_1
XFILLER_138_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[7\].VALID\[6\].TOBUF OVHB\[7\].VALID\[6\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_12362_ _13943_/X VGND VGND VPWR VPWR _12362_/Y sky130_fd_sc_hd__inv_2
XOVHB\[30\].INV _13978_/X VGND VGND VPWR VPWR OVHB\[30\].INV/Y sky130_fd_sc_hd__inv_2
X_11313_ _11343_/CLK line[96] VGND VGND VPWR VPWR _11313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12293_ _12311_/CLK line[32] VGND VGND VPWR VPWR _12293_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11201__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11244_ _11243_/Q _11277_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09456__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11175_ _11191_/CLK line[42] VGND VGND VPWR VPWR _11175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09606__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10126_ _10125_/Q _10157_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13128__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10057_ _10073_/CLK line[43] VGND VGND VPWR VPWR _10057_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06030__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13816_ _13822_/CLK line[83] VGND VGND VPWR VPWR _13816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[2\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _11310_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10487__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13747_ _13747_/A _13762_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10959_ _10958_/Q _10962_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_13678_ _13682_/CLK line[20] VGND VGND VPWR VPWR _13678_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13798__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12629_ _12628_/Q _12642_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07796__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06150_ _06149_/Q _06167_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_05101_ _05093_/CLK line[67] VGND VGND VPWR VPWR _05101_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[13\].TOBUF OVHB\[31\].VALID\[13\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_06081_ _06077_/CLK line[3] VGND VGND VPWR VPWR _06081_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11111__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05032_ _05032_/A _05047_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06205__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10950__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09840_ _09840_/CLK _09841_/X VGND VGND VPWR VPWR _09834_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_99_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08420__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[14\].VALID\[1\].TOBUF OVHB\[14\].VALID\[1\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_09771_ _09912_/A wr VGND VGND VPWR VPWR _09771_/X sky130_fd_sc_hd__and2_1
XFILLER_6_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06983_ _07001_/CLK line[46] VGND VGND VPWR VPWR _06983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13038__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08722_ _13922_/X VGND VGND VPWR VPWR _08722_/Y sky130_fd_sc_hd__inv_2
X_05934_ _05933_/Q _05957_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[13\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07036__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[24\].VALID\[13\].FF OVHB\[24\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[24\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08653_ _08663_/CLK line[32] VGND VGND VPWR VPWR _08653_/Q sky130_fd_sc_hd__dfxtp_1
X_05865_ _05871_/CLK line[47] VGND VGND VPWR VPWR _05865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12877__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07604_ _07603_/Q _07637_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11136__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05796_ _05796_/A _05817_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_08584_ _08583_/Q _08617_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[12\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07535_ _07539_/CLK line[42] VGND VGND VPWR VPWR _07535_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07466_ _07465_/Q _07497_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[0\].FF OVHB\[26\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[26\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06417_ _06421_/CLK line[43] VGND VGND VPWR VPWR _06417_/Q sky130_fd_sc_hd__dfxtp_1
X_09205_ _09204_/Q _09212_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _08125_/CLK sky130_fd_sc_hd__clkbuf_4
X_07397_ _07393_/CLK line[107] VGND VGND VPWR VPWR _07397_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13501__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ _09116_/CLK line[120] VGND VGND VPWR VPWR _09136_/Q sky130_fd_sc_hd__dfxtp_1
X_06348_ _06348_/A _06377_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
X_09067_ _09067_/A _09072_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06279_ _06285_/CLK line[108] VGND VGND VPWR VPWR _06279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08018_ _08000_/CLK line[121] VGND VGND VPWR VPWR _08018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10860__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[5\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09969_ _09968_/Q _09982_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_12980_ _12962_/CLK line[85] VGND VGND VPWR VPWR _12980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[31\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[31\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _11695_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11931_ _11930_/Q _11942_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12787__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11691__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06785__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11862_ _11846_/CLK line[86] VGND VGND VPWR VPWR _11862_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[21\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _08825_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09161__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13601_ _13600_/Q _13622_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_10813_ _10812_/Q _10822_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_11793_ _11793_/A _11802_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[0\].TOBUF OVHB\[20\].VALID\[0\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10100__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13532_ _13528_/CLK line[81] VGND VGND VPWR VPWR _13533_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10744_ _10728_/CLK line[87] VGND VGND VPWR VPWR _10744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13463_ _13463_/A _13482_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_10675_ _10674_/Q _10682_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12414_ _12414_/CLK line[82] VGND VGND VPWR VPWR _12415_/A sky130_fd_sc_hd__dfxtp_1
X_13394_ _13394_/CLK line[18] VGND VGND VPWR VPWR _13394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12027__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12345_ _12344_/Q _12362_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[24\].VALID\[2\].FF OVHB\[24\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[24\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12276_ _12268_/CLK line[19] VGND VGND VPWR VPWR _12276_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11866__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11227_ _11227_/A _11242_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09336__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11158_ _11148_/CLK line[20] VGND VGND VPWR VPWR _11158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10109_ _10109_/A _10122_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_11089_ _11089_/A _11102_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[8\]_A1 _10922_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06695__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05650_ _05650_/A _05677_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[16\]_A0 _10859_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05581_ _05575_/CLK line[45] VGND VGND VPWR VPWR _05581_/Q sky130_fd_sc_hd__dfxtp_1
X_07320_ _07320_/CLK _07321_/X VGND VGND VPWR VPWR _07292_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[20\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _08440_/CLK sky130_fd_sc_hd__clkbuf_4
X_07251_ _13918_/X wr VGND VGND VPWR VPWR _07251_/X sky130_fd_sc_hd__and2_1
XOVHB\[12\].VALID\[6\].TOBUF OVHB\[12\].VALID\[6\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_06202_ _06272_/A VGND VGND VPWR VPWR _06202_/Y sky130_fd_sc_hd__inv_2
XANTENNA__04943__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07182_ _07111_/A VGND VGND VPWR VPWR _07182_/Y sky130_fd_sc_hd__inv_2
X_06133_ _06147_/CLK line[32] VGND VGND VPWR VPWR _06133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[5\].VALID\[10\].TOBUF OVHB\[5\].VALID\[10\].FF/Q OVHB\[5\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_06064_ _06063_/Q _06097_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11776__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[31\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05015_ _05041_/CLK line[42] VGND VGND VPWR VPWR _05015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05774__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09823_ _09822_/Q _09842_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08150__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09754_ _09760_/CLK line[18] VGND VGND VPWR VPWR _09754_/Q sky130_fd_sc_hd__dfxtp_1
X_06966_ _06960_/CLK line[24] VGND VGND VPWR VPWR _06966_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[4\].FF OVHB\[22\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[22\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08705_ _08704_/Q _08722_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_05917_ _05917_/A _05922_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_09685_ _09684_/Q _09702_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_06897_ _06896_/Q _06902_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12400__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08636_ _08646_/CLK line[19] VGND VGND VPWR VPWR _08636_/Q sky130_fd_sc_hd__dfxtp_1
X_05848_ _05836_/CLK line[25] VGND VGND VPWR VPWR _05848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[0\].INV _13983_/Y VGND VGND VPWR VPWR OVHB\[0\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_39_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08567_ _08566_/Q _08582_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11016__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05779_ _05778_/Q _05782_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[7\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07518_ _07518_/CLK line[20] VGND VGND VPWR VPWR _07518_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ _08480_/CLK line[84] VGND VGND VPWR VPWR _08498_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07449_ _07448_/Q _07462_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13231__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05949__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08325__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10460_ _10466_/CLK line[85] VGND VGND VPWR VPWR _10461_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[10\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09119_ _09118_/Q _09142_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
X_10391_ _10390_/Q _10402_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12130_ _12130_/CLK line[95] VGND VGND VPWR VPWR _12131_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10590__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _12061_/A _12082_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[11\].FF OVHB\[20\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[20\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05684__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11012_ _11002_/CLK line[81] VGND VGND VPWR VPWR _11012_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08060__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12963_ _12963_/A _12992_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13406__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11914_ _11934_/CLK line[124] VGND VGND VPWR VPWR _11914_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[3\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12894_ _12902_/CLK line[60] VGND VGND VPWR VPWR _12894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11845_ _11844_/Q _11872_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[6\].FF OVHB\[20\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[20\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11776_ _11776_/CLK line[61] VGND VGND VPWR VPWR _11776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05502__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10765__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13515_ _13515_/CLK _13516_/X VGND VGND VPWR VPWR _13497_/CLK sky130_fd_sc_hd__dlclkp_1
X_10727_ _10726_/Q _10752_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13141__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05859__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[13\].FF OVHB\[10\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[10\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05221__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08235__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13446_ _13552_/A wr VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__and2_1
X_10658_ _10656_/CLK line[62] VGND VGND VPWR VPWR _10659_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12980__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13377_ _13552_/A VGND VGND VPWR VPWR _13377_/Y sky130_fd_sc_hd__inv_2
X_10589_ _10588_/Q _10612_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_12328_ _12352_/CLK line[48] VGND VGND VPWR VPWR _12328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12259_ _12259_/A _12292_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09066__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[12\].TOBUF OVHB\[28\].VALID\[12\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06820_ _06802_/CLK line[85] VGND VGND VPWR VPWR _06820_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13166__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10005__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06751_ _06750_/Q _06762_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13316__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05702_ _05708_/CLK line[86] VGND VGND VPWR VPWR _05703_/A sky130_fd_sc_hd__dfxtp_1
X_09470_ _09482_/CLK line[31] VGND VGND VPWR VPWR _09470_/Q sky130_fd_sc_hd__dfxtp_1
X_06682_ _06682_/CLK line[22] VGND VGND VPWR VPWR _06682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07314__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08421_ _08420_/Q _08442_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[19\].VALID\[7\].FF OVHB\[19\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[19\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05633_ _05633_/A _05642_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08352_ _08358_/CLK line[17] VGND VGND VPWR VPWR _08352_/Q sky130_fd_sc_hd__dfxtp_1
X_05564_ _05568_/CLK line[23] VGND VGND VPWR VPWR _05564_/Q sky130_fd_sc_hd__dfxtp_1
X_07303_ _07302_/Q _07322_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_05495_ _05495_/A _05502_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_08283_ _08282_/Q _08302_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[0\].TOBUF OVHB\[27\].VALID\[0\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_07234_ _07232_/CLK line[18] VGND VGND VPWR VPWR _07235_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13986__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[11\].TOBUF OVHB\[21\].VALID\[11\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12890__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07165_ _07165_/A _07182_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06116_ _06108_/CLK line[19] VGND VGND VPWR VPWR _06116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07096_ _07098_/CLK line[83] VGND VGND VPWR VPWR _07096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[1\].CGAND_A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06047_ _06046_/Q _06062_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09806_ _09912_/A wr VGND VGND VPWR VPWR _09806_/X sky130_fd_sc_hd__and2_1
XFILLER_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07998_ _08000_/CLK line[126] VGND VGND VPWR VPWR _07998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09737_ _09912_/A VGND VGND VPWR VPWR _09737_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06949_ _06948_/Q _06972_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12130__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09668_ _09694_/CLK line[112] VGND VGND VPWR VPWR _09668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07224__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08619_ _08618_/Q _08652_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09598_/Q _09632_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11636_/CLK line[122] VGND VGND VPWR VPWR _11630_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _11561_/A _11592_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13300_/A _13307_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10512_ _10520_/CLK line[123] VGND VGND VPWR VPWR _10512_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _11500_/CLK line[59] VGND VGND VPWR VPWR _11492_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[9\].FF OVHB\[17\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[17\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13896__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13231_ _13213_/CLK line[72] VGND VGND VPWR VPWR _13231_/Q sky130_fd_sc_hd__dfxtp_1
X_10443_ _10442_/Q _10472_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[6\].TOBUF OVHB\[19\].VALID\[6\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ _13161_/Q _13167_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_10374_ _10384_/CLK line[60] VGND VGND VPWR VPWR _10374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12113_ _12109_/CLK line[73] VGND VGND VPWR VPWR _12113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12305__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13093_ _13075_/CLK line[9] VGND VGND VPWR VPWR _13093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05992__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06303__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12044_ _12043_/Q _12047_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09614__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ _12946_/A _12957_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09911__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12877_ _12881_/CLK line[38] VGND VGND VPWR VPWR _12877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06973__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[21\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ _11828_/A _11837_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[13\]_A3 _13562_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10495__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11759_ _11757_/CLK line[39] VGND VGND VPWR VPWR _11759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05589__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05280_ _05278_/CLK line[21] VGND VGND VPWR VPWR _05280_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05886__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13429_ _13439_/CLK line[34] VGND VGND VPWR VPWR _13429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08970_ _08972_/CLK line[58] VGND VGND VPWR VPWR _08970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[13\].FF OVHB\[29\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[29\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06213__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07921_ _07920_/Q _07952_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[0\].VALID\[2\].TOBUF OVHB\[0\].VALID\[2\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_60_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07852_ _07854_/CLK line[59] VGND VGND VPWR VPWR _07852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[25\].VALID\[5\].TOBUF OVHB\[25\].VALID\[5\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_06803_ _06803_/A _06832_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04916__A2 _04918_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07783_ _07782_/Q _07812_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13046__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04995_ _04994_/Q _05012_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
X_09522_ _09521_/Q _09527_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].CG clk OVHB\[31\].CGAND/X VGND VGND VPWR VPWR OVHB\[31\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_06734_ _06740_/CLK line[60] VGND VGND VPWR VPWR _06734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[3\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ _09427_/CLK line[9] VGND VGND VPWR VPWR _09453_/Q sky130_fd_sc_hd__dfxtp_1
X_06665_ _06664_/Q _06692_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07979__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ _08403_/Q _08407_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_05616_ _05632_/CLK line[61] VGND VGND VPWR VPWR _05616_/Q sky130_fd_sc_hd__dfxtp_1
X_09384_ _09383_/Q _09387_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_06596_ _06596_/CLK line[125] VGND VGND VPWR VPWR _06597_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08335_ _08335_/CLK _08336_/X VGND VGND VPWR VPWR _08329_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[3\].CG clk OVHB\[3\].CGAND/X VGND VGND VPWR VPWR OVHB\[3\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_05547_ _05546_/Q _05572_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08266_ _13940_/X wr VGND VGND VPWR VPWR _08266_/X sky130_fd_sc_hd__and2_1
X_05478_ _05476_/CLK line[126] VGND VGND VPWR VPWR _05478_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07217_ _13918_/X VGND VGND VPWR VPWR _07217_/Y sky130_fd_sc_hd__inv_2
X_08197_ _13940_/X VGND VGND VPWR VPWR _08197_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08603__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07148_ _07170_/CLK line[112] VGND VGND VPWR VPWR _07148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07079_ _07079_/A _07112_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10090_ _10100_/CLK line[58] VGND VGND VPWR VPWR _10090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05962__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12800_ _12799_/Q _12817_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_13780_ _13779_/Q _13797_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10992_ _10991_/Q _10997_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07532__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12731_ _12741_/CLK line[99] VGND VGND VPWR VPWR _12731_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12795__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07889__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06793__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07251__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12662_ _12661_/Q _12677_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11605_/CLK line[100] VGND VGND VPWR VPWR _11613_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[4\].TOBUF OVHB\[31\].VALID\[4\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12601_/CLK line[36] VGND VGND VPWR VPWR _12594_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _11543_/Q _11557_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05202__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11475_ _11479_/CLK line[37] VGND VGND VPWR VPWR _11475_/Q sky130_fd_sc_hd__dfxtp_1
X_13214_ _13213_/Q _13237_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08513__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10426_ _10425_/Q _10437_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[22\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12035__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13145_ _13163_/CLK line[47] VGND VGND VPWR VPWR _13145_/Q sky130_fd_sc_hd__dfxtp_1
X_10357_ _10341_/CLK line[38] VGND VGND VPWR VPWR _10357_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07129__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07707__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ _13076_/A _13097_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_10288_ _10288_/A _10297_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_12027_ _12019_/CLK line[33] VGND VGND VPWR VPWR _12027_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07426__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06968__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09344__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13978_ _13979_/A _13979_/B _13979_/C _13979_/D VGND VGND VPWR VPWR _13978_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12929_ _12937_/CLK line[76] VGND VGND VPWR VPWR _12929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06450_ _06464_/CLK line[58] VGND VGND VPWR VPWR _06450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[1\].VALID\[13\].FF OVHB\[1\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[1\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05401_ _05400_/Q _05432_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_06381_ _06380_/Q _06412_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_08120_ _08119_/Q _08127_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_05332_ _05332_/CLK line[59] VGND VGND VPWR VPWR _05332_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04934__A1_N A_h[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08051_ _08033_/CLK line[8] VGND VGND VPWR VPWR _08052_/A sky130_fd_sc_hd__dfxtp_1
X_05263_ _05262_/Q _05292_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09519__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07002_ _07002_/A _07007_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04951__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05194_ _05214_/CLK line[124] VGND VGND VPWR VPWR _05194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[18\].VALID\[10\].TOBUF OVHB\[18\].VALID\[10\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_08953_ _08947_/CLK line[36] VGND VGND VPWR VPWR _08953_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11784__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[4\].FF OVHB\[8\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[8\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07904_ _07903_/Q _07917_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06878__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08884_ _08883_/Q _08897_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09254__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07835_ _07837_/CLK line[37] VGND VGND VPWR VPWR _07835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07766_ _07765_/Q _07777_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04976__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04978_ _05000_/CLK line[16] VGND VGND VPWR VPWR _04978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ _09507_/CLK line[47] VGND VGND VPWR VPWR _09505_/Q sky130_fd_sc_hd__dfxtp_1
X_06717_ _06711_/CLK line[38] VGND VGND VPWR VPWR _06718_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07697_ _07679_/CLK line[102] VGND VGND VPWR VPWR _07697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _09435_/Q _09457_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_06648_ _06647_/Q _06657_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07502__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _09365_/CLK line[97] VGND VGND VPWR VPWR _09367_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11024__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06579_ _06565_/CLK line[103] VGND VGND VPWR VPWR _06579_/Q sky130_fd_sc_hd__dfxtp_1
X_08318_ _08317_/Q _08337_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06118__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ _09297_/Q _09317_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11959__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[11\].FF OVHB\[25\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[25\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08249_ _08257_/CLK line[98] VGND VGND VPWR VPWR _08249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09429__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[3\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08333__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11260_ _11260_/A _11277_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].CGAND _12712_/A wr VGND VGND VPWR VPWR OVHB\[5\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_10_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10211_ _10217_/CLK line[99] VGND VGND VPWR VPWR _10212_/A sky130_fd_sc_hd__dfxtp_1
X_11191_ _11191_/CLK line[35] VGND VGND VPWR VPWR _11191_/Q sky130_fd_sc_hd__dfxtp_1
X_10142_ _10141_/Q _10157_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_10073_ _10073_/CLK line[36] VGND VGND VPWR VPWR _10074_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05692__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05047__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13901_ _13907_/X wr VGND VGND VPWR VPWR _13901_/X sky130_fd_sc_hd__and2_1
XOVHB\[7\].VALID\[2\].TOBUF OVHB\[7\].VALID\[2\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_13832_ _13907_/X VGND VGND VPWR VPWR _13832_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13763_ _13763_/CLK line[64] VGND VGND VPWR VPWR _13763_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[13\].FF OVHB\[15\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[15\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[6\].FF OVHB\[6\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[6\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10975_ _10977_/CLK line[79] VGND VGND VPWR VPWR _10976_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _12713_/Q _12747_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08508__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13694_ _13693_/Q _13727_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _12667_/CLK line[74] VGND VGND VPWR VPWR _12645_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06028__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12576_ _12576_/A _12607_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10773__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11535_/CLK line[75] VGND VGND VPWR VPWR _11527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05867__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08243__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11458_ _11457_/Q _11487_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_10409_ _10405_/CLK line[76] VGND VGND VPWR VPWR _10409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11389_ _11395_/CLK line[12] VGND VGND VPWR VPWR _11390_/A sky130_fd_sc_hd__dfxtp_1
X_13128_ _13120_/CLK line[25] VGND VGND VPWR VPWR _13128_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06341__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05950_ _05950_/A _05957_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_13059_ _13059_/A _13062_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[20\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05881_ _05871_/CLK line[40] VGND VGND VPWR VPWR _05882_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11109__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07620_ _07619_/Q _07637_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10013__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05107__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07551_ _07539_/CLK line[35] VGND VGND VPWR VPWR _07552_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10948__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13324__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13902__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06502_ _06501_/Q _06517_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08418__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07482_ _07481_/Q _07497_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_09221_ _09241_/CLK line[45] VGND VGND VPWR VPWR _09222_/A sky130_fd_sc_hd__dfxtp_1
X_06433_ _06421_/CLK line[36] VGND VGND VPWR VPWR _06433_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13621__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09152_ _09151_/Q _09177_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06364_ _06363_/Q _06377_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06516__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08103_ _08113_/CLK line[46] VGND VGND VPWR VPWR _08104_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[8\].FF OVHB\[4\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[4\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05315_ _05299_/CLK line[37] VGND VGND VPWR VPWR _05315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10683__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06295_ _06285_/CLK line[101] VGND VGND VPWR VPWR _06296_/A sky130_fd_sc_hd__dfxtp_1
X_09083_ _09085_/CLK line[110] VGND VGND VPWR VPWR _09084_/A sky130_fd_sc_hd__dfxtp_1
X_08034_ _08033_/Q _08057_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_05246_ _05246_/A _05257_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[26\]_A2 _06521_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05177_ _05157_/CLK line[102] VGND VGND VPWR VPWR _05177_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07992__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09985_ _10011_/CLK line[10] VGND VGND VPWR VPWR _09985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08936_ _08935_/Q _08967_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09562__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08867_ _08869_/CLK line[11] VGND VGND VPWR VPWR _08867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07818_ _07817_/Q _07847_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09281__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _08798_/A _08827_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05017__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10858__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07749_ _07773_/CLK line[12] VGND VGND VPWR VPWR _07749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10760_ _10759_/Q _10787_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07232__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09419_ _09418_/Q _09422_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_10691_ _10707_/CLK line[77] VGND VGND VPWR VPWR _10691_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ _12430_/CLK _12431_/X VGND VGND VPWR VPWR _12414_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11689__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12361_ _13943_/X wr VGND VGND VPWR VPWR _12361_/X sky130_fd_sc_hd__and2_1
XANTENNA__09159__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[7\].TOBUF OVHB\[5\].VALID\[7\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_11312_ _11311_/A VGND VGND VPWR VPWR _11312_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09737__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12292_ _13943_/X VGND VGND VPWR VPWR _12292_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11243_ _11251_/CLK line[64] VGND VGND VPWR VPWR _11243_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08998__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09456__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11174_ _11173_/Q _11207_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12313__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10125_ _10145_/CLK line[74] VGND VGND VPWR VPWR _10125_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[19\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07407__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10056_ _10055_/Q _10087_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09622__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13815_ _13814_/Q _13832_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13746_ _13746_/CLK line[51] VGND VGND VPWR VPWR _13747_/A sky130_fd_sc_hd__dfxtp_1
X_10958_ _10930_/CLK line[57] VGND VGND VPWR VPWR _10958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13677_ _13676_/Q _13692_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_10889_ _10889_/A _10892_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11242__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ _12638_/CLK line[52] VGND VGND VPWR VPWR _12628_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06981__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12559_ _12558_/Q _12572_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05597__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05100_ _05099_/Q _05117_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_06080_ _06079_/Q _06097_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[0\].FF OVHB\[13\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[13\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05031_ _05041_/CLK line[35] VGND VGND VPWR VPWR _05032_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[4\].FF OVHB\[30\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[30\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12223__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09770_ _09770_/CLK _09771_/X VGND VGND VPWR VPWR _09760_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[11\].VALID\[11\].FF OVHB\[11\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[11\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06982_ _06982_/A _07007_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08721_ _13922_/X wr VGND VGND VPWR VPWR _08721_/X sky130_fd_sc_hd__and2_1
XANTENNA__06221__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[2\].TOBUF OVHB\[12\].VALID\[2\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_05933_ _05929_/CLK line[78] VGND VGND VPWR VPWR _05933_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11417__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _13922_/X VGND VGND VPWR VPWR _08652_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05864_ _05864_/A _05887_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09532__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07603_ _07633_/CLK line[64] VGND VGND VPWR VPWR _07603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10678__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11136__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08583_ _08609_/CLK line[0] VGND VGND VPWR VPWR _08583_/Q sky130_fd_sc_hd__dfxtp_1
X_05795_ _05799_/CLK line[15] VGND VGND VPWR VPWR _05796_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13054__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07534_ _07533_/Q _07567_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08148__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13989__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07465_ _07467_/CLK line[10] VGND VGND VPWR VPWR _07465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09204_ _09200_/CLK line[23] VGND VGND VPWR VPWR _09204_/Q sky130_fd_sc_hd__dfxtp_1
X_06416_ _06415_/Q _06447_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
X_07396_ _07395_/Q _07427_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09135_ _09134_/Q _09142_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_06347_ _06353_/CLK line[11] VGND VGND VPWR VPWR _06348_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11302__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09066_ _09068_/CLK line[88] VGND VGND VPWR VPWR _09067_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[5\].FF OVHB\[29\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[29\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06278_ _06277_/Q _06307_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08017_ _08016_/Q _08022_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05229_ _05253_/CLK line[12] VGND VGND VPWR VPWR _05229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09707__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07077__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08611__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13229__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09968_ _09978_/CLK line[116] VGND VGND VPWR VPWR _09968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[11\].VALID\[2\].FF OVHB\[11\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[11\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12711__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08919_ _08919_/A _08932_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09899_ _09898_/Q _09912_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11930_ _11934_/CLK line[117] VGND VGND VPWR VPWR _11930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05970__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10588__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11861_ _11861_/A _11872_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13600_ _13598_/CLK line[127] VGND VGND VPWR VPWR _13600_/Q sky130_fd_sc_hd__dfxtp_1
X_10812_ _10804_/CLK line[118] VGND VGND VPWR VPWR _10812_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08058__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11792_ _11776_/CLK line[54] VGND VGND VPWR VPWR _11793_/A sky130_fd_sc_hd__dfxtp_1
X_13531_ _13530_/Q _13552_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_10743_ _10743_/A _10752_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DECH.DEC0.AND1_B A_h[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07897__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13462_ _13468_/CLK line[49] VGND VGND VPWR VPWR _13463_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10674_ _10656_/CLK line[55] VGND VGND VPWR VPWR _10674_/Q sky130_fd_sc_hd__dfxtp_1
X_12413_ _12413_/A _12432_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_13393_ _13392_/Q _13412_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11212__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12344_ _12352_/CLK line[50] VGND VGND VPWR VPWR _12344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08371__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05210__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[12\].TOBUF OVHB\[8\].VALID\[12\].FF/Q OVHB\[8\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_12275_ _12274_/Q _12292_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11226_ _11216_/CLK line[51] VGND VGND VPWR VPWR _11227_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08521__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13139__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12043__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11157_ _11156_/Q _11172_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07137__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[7\].FF OVHB\[27\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[27\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10108_ _10100_/CLK line[52] VGND VGND VPWR VPWR _10109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12978__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11088_ _11090_/CLK line[116] VGND VGND VPWR VPWR _11089_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[13\].FF OVHB\[6\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[6\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[8\]_A2 _10992_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10039_ _10038_/Q _10052_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[17\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05580_ _05579_/Q _05607_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[16\]_A1 _07009_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08546__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13729_ _13729_/A _13762_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13602__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[11\].TOBUF OVHB\[1\].VALID\[11\].FF/Q OVHB\[1\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_07250_ _07250_/CLK _07251_/X VGND VGND VPWR VPWR _07232_/CLK sky130_fd_sc_hd__dlclkp_1
X_06201_ _06272_/A wr VGND VGND VPWR VPWR _06201_/X sky130_fd_sc_hd__and2_1
XANTENNA__12218__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07181_ _07111_/A wr VGND VGND VPWR VPWR _07181_/X sky130_fd_sc_hd__and2_1
XOVHB\[10\].VALID\[7\].TOBUF OVHB\[10\].VALID\[7\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06132_ _06272_/A VGND VGND VPWR VPWR _06132_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05120__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[19\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _07810_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_117_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06063_ _06077_/CLK line[0] VGND VGND VPWR VPWR _06063_/Q sky130_fd_sc_hd__dfxtp_1
X_05014_ _05013_/Q _05047_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09822_ _09834_/CLK line[49] VGND VGND VPWR VPWR _09822_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07047__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12888__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09753_ _09753_/A _09772_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_06965_ _06964_/Q _06972_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11792__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08704_ _08710_/CLK line[50] VGND VGND VPWR VPWR _08704_/Q sky130_fd_sc_hd__dfxtp_1
X_05916_ _05902_/CLK line[56] VGND VGND VPWR VPWR _05917_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06886__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09684_ _09694_/CLK line[114] VGND VGND VPWR VPWR _09684_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10051__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09262__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06896_ _06892_/CLK line[120] VGND VGND VPWR VPWR _06896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08635_ _08634_/Q _08652_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05847_ _05846_/Q _05852_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10201__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08566_ _08560_/CLK line[115] VGND VGND VPWR VPWR _08566_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[9\].FF OVHB\[25\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[25\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05778_ _05756_/CLK line[121] VGND VGND VPWR VPWR _05778_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ _07516_/Q _07532_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _08496_/Q _08512_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07448_ _07446_/CLK line[116] VGND VGND VPWR VPWR _07448_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07510__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12128__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07379_ _07378_/Q _07392_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_09118_ _09116_/CLK line[126] VGND VGND VPWR VPWR _09118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06126__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10390_ _10384_/CLK line[53] VGND VGND VPWR VPWR _10390_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11967__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09049_ _09048_/Q _09072_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10226__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09437__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ _12072_/CLK line[63] VGND VGND VPWR VPWR _12061_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11011_ _11010_/Q _11032_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04937__B1 A_h[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12962_ _12962_/CLK line[91] VGND VGND VPWR VPWR _12963_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11913_ _11913_/A _11942_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VALID\[2\].TOBUF OVHB\[19\].VALID\[2\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_12893_ _12892_/Q _12922_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13272__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11844_ _11846_/CLK line[92] VGND VGND VPWR VPWR _11844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09900__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11775_ _11774_/Q _11802_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13514_ _13513_/Q _13517_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_10726_ _10728_/CLK line[93] VGND VGND VPWR VPWR _10726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13445_ _13445_/CLK _13446_/X VGND VGND VPWR VPWR _13439_/CLK sky130_fd_sc_hd__dlclkp_1
X_10657_ _10657_/A _10682_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[24\].VALID\[13\].TOBUF OVHB\[24\].VALID\[13\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06036__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13376_ _13552_/A wr VGND VGND VPWR VPWR _13376_/X sky130_fd_sc_hd__and2_1
X_10588_ _10594_/CLK line[30] VGND VGND VPWR VPWR _10588_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11877__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10781__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12327_ _13943_/X VGND VGND VPWR VPWR _12327_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05875__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08251__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12258_ _12268_/CLK line[16] VGND VGND VPWR VPWR _12259_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[30\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11209_ _11208_/Q _11242_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13447__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12189_ _12188_/Q _12222_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13166__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04928__B1 A_h[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06750_ _06740_/CLK line[53] VGND VGND VPWR VPWR _06750_/Q sky130_fd_sc_hd__dfxtp_1
X_05701_ _05701_/A _05712_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_06681_ _06681_/A _06692_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11117__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08420_ _08410_/CLK line[63] VGND VGND VPWR VPWR _08420_/Q sky130_fd_sc_hd__dfxtp_1
X_05632_ _05632_/CLK line[54] VGND VGND VPWR VPWR _05633_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09810__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10956__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08351_ _08351_/A _08372_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_05563_ _05562_/Q _05572_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13332__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07302_ _07292_/CLK line[49] VGND VGND VPWR VPWR _07302_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08426__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08282_ _08282_/CLK line[113] VGND VGND VPWR VPWR _08282_/Q sky130_fd_sc_hd__dfxtp_1
X_05494_ _05476_/CLK line[119] VGND VGND VPWR VPWR _05495_/A sky130_fd_sc_hd__dfxtp_1
X_07233_ _07232_/Q _07252_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[1\].TOBUF OVHB\[25\].VALID\[1\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_118_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07164_ _07170_/CLK line[114] VGND VGND VPWR VPWR _07165_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10691__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06115_ _06114_/Q _06132_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
X_07095_ _07094_/Q _07112_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05785__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06046_ _06050_/CLK line[115] VGND VGND VPWR VPWR _06046_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].CGAND_A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[11\].FF OVHB\[2\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[2\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[5\].CGAND_A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09805_ _09805_/CLK _09806_/X VGND VGND VPWR VPWR _09793_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__04919__B1 A_h[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07997_ _07997_/A _08022_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13507__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09736_ _09912_/A wr VGND VGND VPWR VPWR _09736_/X sky130_fd_sc_hd__and2_1
X_06948_ _06960_/CLK line[30] VGND VGND VPWR VPWR _06948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09667_ _09632_/A VGND VGND VPWR VPWR _09667_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06879_ _06879_/A _06902_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08618_ _08646_/CLK line[16] VGND VGND VPWR VPWR _08618_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09626_/CLK line[80] VGND VGND VPWR VPWR _09598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05025__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08548_/Q _08582_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10866__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13242__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11588_/CLK line[90] VGND VGND VPWR VPWR _11561_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07240__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[30\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ _10511_/A _10542_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _11490_/Q _11522_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13229_/Q _13237_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10442_ _10466_/CLK line[91] VGND VGND VPWR VPWR _10442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13161_ _13163_/CLK line[40] VGND VGND VPWR VPWR _13161_/Q sky130_fd_sc_hd__dfxtp_1
X_10373_ _10372_/Q _10402_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[7\].TOBUF OVHB\[17\].VALID\[7\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09167__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12112_ _12111_/Q _12117_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13092_ _13091_/Q _13097_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_12043_ _12019_/CLK line[41] VGND VGND VPWR VPWR _12043_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10106__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[31\].VALID\[0\].TOBUF OVHB\[31\].VALID\[0\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_46_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13417__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12321__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07415__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12945_ _12937_/CLK line[69] VGND VGND VPWR VPWR _12946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12876_ _12875_/Q _12887_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[21\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11827_ _11823_/CLK line[70] VGND VGND VPWR VPWR _11828_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XMUX.MUX\[0\] _06904_/Z _10894_/Z _05084_/Z _13554_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[0] sky130_fd_sc_hd__mux4_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11758_ _11757_/Q _11767_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07150__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10709_ _10707_/CLK line[71] VGND VGND VPWR VPWR _10709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11689_ _11691_/CLK line[7] VGND VGND VPWR VPWR _11690_/A sky130_fd_sc_hd__dfxtp_1
X_13428_ _13427_/Q _13447_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[11\].FF OVHB\[16\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[16\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13359_ _13347_/CLK line[2] VGND VGND VPWR VPWR _13360_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09077__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ _07946_/CLK line[90] VGND VGND VPWR VPWR _07920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12081__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[19\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07851_ _07850_/Q _07882_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06802_ _06802_/CLK line[91] VGND VGND VPWR VPWR _06803_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12231__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04949__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13905__A A[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07782_ _07788_/CLK line[27] VGND VGND VPWR VPWR _07782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04994_ _05000_/CLK line[18] VGND VGND VPWR VPWR _04994_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[6\].TOBUF OVHB\[23\].VALID\[6\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__07325__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09521_ _09507_/CLK line[40] VGND VGND VPWR VPWR _09521_/Q sky130_fd_sc_hd__dfxtp_1
X_06733_ _06732_/Q _06762_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _09451_/Q _09457_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_06664_ _06682_/CLK line[28] VGND VGND VPWR VPWR _06664_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09540__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08403_ _08383_/CLK line[41] VGND VGND VPWR VPWR _08403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05615_ _05614_/Q _05642_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_09383_ _09365_/CLK line[105] VGND VGND VPWR VPWR _09383_/Q sky130_fd_sc_hd__dfxtp_1
X_06595_ _06594_/Q _06622_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[29\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08334_ _08333_/Q _08337_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08156__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05546_ _05568_/CLK line[29] VGND VGND VPWR VPWR _05546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ _08265_/CLK _08266_/X VGND VGND VPWR VPWR _08257_/CLK sky130_fd_sc_hd__dlclkp_1
X_05477_ _05476_/Q _05502_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12256__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07216_ _13918_/X wr VGND VGND VPWR VPWR _07216_/X sky130_fd_sc_hd__and2_1
X_08196_ _13940_/X wr VGND VGND VPWR VPWR _08196_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.MUX\[29\]_A0 _10867_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07147_ _07111_/A VGND VGND VPWR VPWR _07147_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12406__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06404__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07078_ _07098_/CLK line[80] VGND VGND VPWR VPWR _07079_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06029_ _06028_/Q _06062_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09715__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09719_ _09721_/CLK line[2] VGND VGND VPWR VPWR _09719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10991_ _10977_/CLK line[72] VGND VGND VPWR VPWR _10991_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11980__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].CGAND _13940_/X wr VGND VGND VPWR VPWR OVHB\[1\].CGAND/X sky130_fd_sc_hd__and2_4
X_12730_ _12729_/Q _12747_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12667_/CLK line[67] VGND VGND VPWR VPWR _12661_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10596__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11611_/Q _11627_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08066__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12592_ _12591_/Q _12607_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _11535_/CLK line[68] VGND VGND VPWR VPWR _11543_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11474_ _11474_/A _11487_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_13213_ _13213_/CLK line[78] VGND VGND VPWR VPWR _13213_/Q sky130_fd_sc_hd__dfxtp_1
X_10425_ _10405_/CLK line[69] VGND VGND VPWR VPWR _10425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11220__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13144_ _13143_/Q _13167_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06314__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10356_ _10355_/Q _10367_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[9\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _13725_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_83_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13075_ _13075_/CLK line[15] VGND VGND VPWR VPWR _13076_/A sky130_fd_sc_hd__dfxtp_1
X_10287_ _10277_/CLK line[6] VGND VGND VPWR VPWR _10288_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12026_ _12025_/Q _12047_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13147__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12986__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ _13979_/B _13979_/A _13979_/C _13979_/D VGND VGND VPWR VPWR _13977_/X sky130_fd_sc_hd__and4b_4
XFILLER_4_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12928_ _12927_/Q _12957_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12859_ _12881_/CLK line[44] VGND VGND VPWR VPWR _12859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05400_ _05424_/CLK line[90] VGND VGND VPWR VPWR _05400_/Q sky130_fd_sc_hd__dfxtp_1
X_06380_ _06408_/CLK line[26] VGND VGND VPWR VPWR _06380_/Q sky130_fd_sc_hd__dfxtp_1
X_05331_ _05330_/Q _05362_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[11\].TOBUF OVHB\[14\].VALID\[11\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _11065_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13610__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08050_ _08049_/Q _08057_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08704__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05262_ _05278_/CLK line[27] VGND VGND VPWR VPWR _05262_/Q sky130_fd_sc_hd__dfxtp_1
X_07001_ _07001_/CLK line[40] VGND VGND VPWR VPWR _07002_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05193_ _05193_/A _05222_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08952_ _08951_/Q _08967_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07903_ _07905_/CLK line[68] VGND VGND VPWR VPWR _07903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08883_ _08869_/CLK line[4] VGND VGND VPWR VPWR _08883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07834_ _07833_/Q _07847_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07055__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12896__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07765_ _07773_/CLK line[5] VGND VGND VPWR VPWR _07765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04977_ _05152_/A VGND VGND VPWR VPWR _04977_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__04976__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06716_ _06715_/Q _06727_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_09504_ _09503_/Q _09527_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06894__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07696_ _07695_/Q _07707_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09270__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09435_ _09427_/CLK line[15] VGND VGND VPWR VPWR _09435_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06647_ _06633_/CLK line[6] VGND VGND VPWR VPWR _06647_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _09366_/A _09387_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06578_ _06577_/Q _06587_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05303__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08317_ _08329_/CLK line[1] VGND VGND VPWR VPWR _08317_/Q sky130_fd_sc_hd__dfxtp_1
X_05529_ _05519_/CLK line[7] VGND VGND VPWR VPWR _05530_/A sky130_fd_sc_hd__dfxtp_1
X_09297_ _09307_/CLK line[65] VGND VGND VPWR VPWR _09297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13520__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _08247_/Q _08267_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12136__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[3\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08179_ _08175_/CLK line[66] VGND VGND VPWR VPWR _08179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10210_ _10210_/A _10227_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[28\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _10680_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11190_ _11189_/Q _11207_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10141_ _10145_/CLK line[67] VGND VGND VPWR VPWR _10141_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[11\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09445__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10072_ _10071_/Q _10087_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13900_ _13900_/CLK _13901_/X VGND VGND VPWR VPWR _13882_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_87_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13831_ _13907_/X wr VGND VGND VPWR VPWR _13831_/X sky130_fd_sc_hd__and2_1
XOVHB\[5\].VALID\[3\].TOBUF OVHB\[5\].VALID\[3\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_29_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[3\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13762_ _13907_/X VGND VGND VPWR VPWR _13762_/Y sky130_fd_sc_hd__inv_2
X_10974_ _10973_/Q _10997_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09180__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _12741_/CLK line[96] VGND VGND VPWR VPWR _12713_/Q sky130_fd_sc_hd__dfxtp_1
X_13693_ _13701_/CLK line[32] VGND VGND VPWR VPWR _13693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[0\].FF OVHB\[21\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[21\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ _12643_/Q _12677_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _12601_/CLK line[42] VGND VGND VPWR VPWR _12576_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[22\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _11525_/Q _11557_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11457_ _11479_/CLK line[43] VGND VGND VPWR VPWR _11457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].CG clk OVHB\[21\].CGAND/X VGND VGND VPWR VPWR OVHB\[21\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_125_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06044__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10408_ _10407_/Q _10437_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_11388_ _11387_/Q _11417_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06622__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11885__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10339_ _10341_/CLK line[44] VGND VGND VPWR VPWR _10339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06979__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[0\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13127_ _13127_/A _13132_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05883__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06341__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09355__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13058_ _13050_/CLK line[121] VGND VGND VPWR VPWR _13059_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[27\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _10295_/CLK sky130_fd_sc_hd__clkbuf_4
X_12009_ _12008_/Q _12012_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
X_05880_ _05879_/Q _05887_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _07425_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07550_ _07549_/Q _07567_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07603__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06501_ _06489_/CLK line[67] VGND VGND VPWR VPWR _06501_/Q sky130_fd_sc_hd__dfxtp_1
X_07481_ _07467_/CLK line[3] VGND VGND VPWR VPWR _07481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11125__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09220_ _09219_/Q _09247_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_06432_ _06431_/Q _06447_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06219__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09151_ _09147_/CLK line[13] VGND VGND VPWR VPWR _09151_/Q sky130_fd_sc_hd__dfxtp_1
X_06363_ _06353_/CLK line[4] VGND VGND VPWR VPWR _06363_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[11\].FF OVHB\[7\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[7\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08102_ _08101_/Q _08127_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06516__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05314_ _05313_/Q _05327_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_09082_ _09081_/Q _09107_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08434__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06294_ _06293_/Q _06307_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_08033_ _08033_/CLK line[14] VGND VGND VPWR VPWR _08033_/Q sky130_fd_sc_hd__dfxtp_1
X_05245_ _05253_/CLK line[5] VGND VGND VPWR VPWR _05246_/A sky130_fd_sc_hd__dfxtp_1
X_05176_ _05175_/Q _05187_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[26\]_A3 _13591_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[5\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05793__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09984_ _09983_/Q _10017_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_08935_ _08947_/CLK line[42] VGND VGND VPWR VPWR _08935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08866_ _08865_/Q _08897_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_07817_ _07837_/CLK line[43] VGND VGND VPWR VPWR _07817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08797_ _08823_/CLK line[107] VGND VGND VPWR VPWR _08798_/A sky130_fd_sc_hd__dfxtp_1
X_07748_ _07747_/Q _07777_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08609__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07679_ _07679_/CLK line[108] VGND VGND VPWR VPWR _07680_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[16\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _07040_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11035__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09418_ _09414_/CLK line[121] VGND VGND VPWR VPWR _09418_/Q sky130_fd_sc_hd__dfxtp_1
X_10690_ _10689_/Q _10717_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05033__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10874__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09349_ _09348_/Q _09352_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13250__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05968__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12360_ _12360_/CLK _12361_/X VGND VGND VPWR VPWR _12352_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08344__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[18\].VALID\[3\].FF OVHB\[18\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[18\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11311_ _11311_/A wr VGND VGND VPWR VPWR _11311_/X sky130_fd_sc_hd__and2_1
X_12291_ _13943_/X wr VGND VGND VPWR VPWR _12291_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[28\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[8\].TOBUF OVHB\[3\].VALID\[8\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_101_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11242_ _11311_/A VGND VGND VPWR VPWR _11242_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11173_ _11191_/CLK line[32] VGND VGND VPWR VPWR _11173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10124_ _10123_/Q _10157_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[25\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10114__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10055_ _10073_/CLK line[42] VGND VGND VPWR VPWR _10055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05208__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04933__A1_N A_h[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13425__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13814_ _13822_/CLK line[82] VGND VGND VPWR VPWR _13814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08519__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07423__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13745_ _13744_/Q _13762_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_10957_ _10956_/Q _10962_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13676_ _13682_/CLK line[19] VGND VGND VPWR VPWR _13676_/Q sky130_fd_sc_hd__dfxtp_1
X_10888_ _10872_/CLK line[25] VGND VGND VPWR VPWR _10889_/A sky130_fd_sc_hd__dfxtp_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _12626_/Q _12642_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[15\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _06655_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12558_ _12560_/CLK line[20] VGND VGND VPWR VPWR _12558_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11509_ _11508_/Q _11522_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12489_ _12488_/Q _12502_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_05030_ _05029_/Q _05047_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09085__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[16\].VALID\[5\].FF OVHB\[16\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[16\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06981_ _07001_/CLK line[45] VGND VGND VPWR VPWR _06982_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08720_ _08720_/CLK _08721_/X VGND VGND VPWR VPWR _08710_/CLK sky130_fd_sc_hd__dlclkp_1
X_05932_ _05931_/Q _05957_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10024__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05118__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[3\].TOBUF OVHB\[10\].VALID\[3\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_08651_ _13922_/X wr VGND VGND VPWR VPWR _08651_/X sky130_fd_sc_hd__and2_1
X_05863_ _05871_/CLK line[46] VGND VGND VPWR VPWR _05864_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07602_ _07672_/A VGND VGND VPWR VPWR _07602_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08582_ _13921_/X VGND VGND VPWR VPWR _08582_/Y sky130_fd_sc_hd__inv_2
XANTENNA__04957__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05794_ _05793_/Q _05817_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07333__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07533_ _07539_/CLK line[32] VGND VGND VPWR VPWR _07533_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07464_ _07463_/Q _07497_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_06415_ _06421_/CLK line[42] VGND VGND VPWR VPWR _06415_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05431__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09203_ _09202_/Q _09212_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_07395_ _07393_/CLK line[106] VGND VGND VPWR VPWR _07395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09134_ _09116_/CLK line[119] VGND VGND VPWR VPWR _09134_/Q sky130_fd_sc_hd__dfxtp_1
X_06346_ _06345_/Q _06377_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09065_ _09064_/Q _09072_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_06277_ _06285_/CLK line[107] VGND VGND VPWR VPWR _06277_/Q sky130_fd_sc_hd__dfxtp_1
X_08016_ _08000_/CLK line[120] VGND VGND VPWR VPWR _08016_/Q sky130_fd_sc_hd__dfxtp_1
X_05228_ _05227_/Q _05257_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12414__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05159_ _05157_/CLK line[108] VGND VGND VPWR VPWR _05159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07508__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09967_ _09966_/Q _09982_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12711__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08918_ _08922_/CLK line[20] VGND VGND VPWR VPWR _08919_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09898_ _09908_/CLK line[84] VGND VGND VPWR VPWR _09898_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09723__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05606__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08849_ _08848_/Q _08862_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_11860_ _11846_/CLK line[85] VGND VGND VPWR VPWR _11861_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[7\].FF OVHB\[14\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[14\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10811_ _10810_/Q _10822_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_11791_ _11790_/Q _11802_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13530_ _13528_/CLK line[95] VGND VGND VPWR VPWR _13530_/Q sky130_fd_sc_hd__dfxtp_1
X_10742_ _10728_/CLK line[86] VGND VGND VPWR VPWR _10743_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[13\].TOBUF OVHB\[4\].VALID\[13\].FF/Q OVHB\[4\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_10673_ _10672_/Q _10682_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_13461_ _13460_/Q _13482_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05698__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08074__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12412_ _12414_/CLK line[81] VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08652__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13392_ _13394_/CLK line[17] VGND VGND VPWR VPWR _13392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _12342_/Q _12362_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08371__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12274_ _12268_/CLK line[18] VGND VGND VPWR VPWR _12274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11225_ _11224_/Q _11242_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06322__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11156_ _11148_/CLK line[19] VGND VGND VPWR VPWR _11156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10107_ _10107_/A _10122_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_11087_ _11086_/Q _11102_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09633__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10779__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10038_ _10042_/CLK line[20] VGND VGND VPWR VPWR _10038_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[8\]_A3 _13582_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13155__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08249__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08827__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[16\]_A2 _05119_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _11988_/Q _12012_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08546__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13728_ _13746_/CLK line[48] VGND VGND VPWR VPWR _13729_/A sky130_fd_sc_hd__dfxtp_1
X_13659_ _13659_/A _13692_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11403__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06200_ _06200_/CLK _06201_/X VGND VGND VPWR VPWR _06186_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[12\].VALID\[9\].FF OVHB\[12\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[12\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07180_ _07180_/CLK _07181_/X VGND VGND VPWR VPWR _07170_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06131_ _06272_/A wr VGND VGND VPWR VPWR _06131_/X sky130_fd_sc_hd__and2_1
XANTENNA__09808__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08712__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06062_ _13910_/X VGND VGND VPWR VPWR _06062_/Y sky130_fd_sc_hd__inv_2
X_05013_ _05041_/CLK line[32] VGND VGND VPWR VPWR _05013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09821_ _09820_/Q _09842_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09752_ _09760_/CLK line[17] VGND VGND VPWR VPWR _09753_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10332__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06964_ _06960_/CLK line[23] VGND VGND VPWR VPWR _06964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08703_ _08703_/A _08722_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_05915_ _05914_/Q _05922_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10689__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06895_ _06894_/Q _06902_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_09683_ _09683_/A _09702_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13065__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10051__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05846_ _05836_/CLK line[24] VGND VGND VPWR VPWR _05846_/Q sky130_fd_sc_hd__dfxtp_1
X_08634_ _08646_/CLK line[18] VGND VGND VPWR VPWR _08634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07063__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08565_ _08564_/Q _08582_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_05777_ _05777_/A _05782_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07998__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ _07518_/CLK line[19] VGND VGND VPWR VPWR _07516_/Q sky130_fd_sc_hd__dfxtp_1
X_08496_ _08480_/CLK line[83] VGND VGND VPWR VPWR _08496_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07447_ _07447_/A _07462_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11313__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[30\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[24\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07378_ _07380_/CLK line[84] VGND VGND VPWR VPWR _07378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05311__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09117_ _09116_/Q _09142_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_06329_ _06328_/Q _06342_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10507__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09048_ _09068_/CLK line[94] VGND VGND VPWR VPWR _09048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08622__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10226__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12144__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07238__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11010_ _11002_/CLK line[95] VGND VGND VPWR VPWR _11010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04937__B2 _04937_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09453__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ _12960_/Q _12992_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11912_ _11934_/CLK line[123] VGND VGND VPWR VPWR _11913_/A sky130_fd_sc_hd__dfxtp_1
X_12892_ _12902_/CLK line[59] VGND VGND VPWR VPWR _12892_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _13340_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[17\].VALID\[3\].TOBUF OVHB\[17\].VALID\[3\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11843_ _11842_/Q _11872_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[0\].FF OVHB\[7\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[7\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13703__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[14\].TOBUF OVHB\[20\].VALID\[14\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[18\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06167__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11774_ _11776_/CLK line[60] VGND VGND VPWR VPWR _11774_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07701__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13513_ _13497_/CLK line[73] VGND VGND VPWR VPWR _13513_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12319__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10725_ _10724_/Q _10752_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11801__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13444_ _13443_/Q _13447_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_10656_ _10656_/CLK line[61] VGND VGND VPWR VPWR _10657_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[22\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13375_ _13375_/CLK _13376_/X VGND VGND VPWR VPWR _13347_/CLK sky130_fd_sc_hd__dlclkp_1
X_10587_ _10586_/Q _10612_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09628__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12326_ _13943_/X wr VGND VGND VPWR VPWR _12326_/X sky130_fd_sc_hd__and2_1
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12054__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12257_ _13943_/X VGND VGND VPWR VPWR _12257_/Y sky130_fd_sc_hd__inv_2
XOVHB\[26\].V OVHB\[26\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[26\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07148__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06052__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11208_ _11216_/CLK line[48] VGND VGND VPWR VPWR _11208_/Q sky130_fd_sc_hd__dfxtp_1
X_12188_ _12204_/CLK line[112] VGND VGND VPWR VPWR _12188_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11893__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06987__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11139_ _11138_/Q _11172_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09363__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05700_ _05708_/CLK line[85] VGND VGND VPWR VPWR _05701_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10302__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06680_ _06682_/CLK line[21] VGND VGND VPWR VPWR _06681_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07461__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05631_ _05630_/Q _05642_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_08350_ _08358_/CLK line[31] VGND VGND VPWR VPWR _08351_/A sky130_fd_sc_hd__dfxtp_1
X_05562_ _05568_/CLK line[22] VGND VGND VPWR VPWR _05562_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07611__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07301_ _07300_/Q _07322_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12229__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08281_ _08280_/Q _08302_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[6\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _12955_/CLK sky130_fd_sc_hd__clkbuf_4
X_05493_ _05493_/A _05502_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11133__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07232_ _07232_/CLK line[17] VGND VGND VPWR VPWR _07232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06227__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[2\].FF OVHB\[5\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[5\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[2\].TOBUF OVHB\[23\].VALID\[2\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_07163_ _07162_/Q _07182_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09538__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06114_ _06108_/CLK line[18] VGND VGND VPWR VPWR _06114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07094_ _07098_/CLK line[82] VGND VGND VPWR VPWR _07094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06045_ _06044_/Q _06062_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].V OVHB\[17\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[17\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07636__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[5\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09804_ _09804_/A _09807_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].CGAND_A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04919__B2 _04919_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07996_ _08000_/CLK line[125] VGND VGND VPWR VPWR _07997_/A sky130_fd_sc_hd__dfxtp_1
X_09735_ _09735_/CLK _09736_/X VGND VGND VPWR VPWR _09721_/CLK sky130_fd_sc_hd__dlclkp_1
X_06947_ _06947_/A _06972_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10997__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11308__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].CGAND_A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09666_ _09632_/A wr VGND VGND VPWR VPWR _09666_/X sky130_fd_sc_hd__and2_1
X_06878_ _06892_/CLK line[126] VGND VGND VPWR VPWR _06879_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _13922_/X VGND VGND VPWR VPWR _08617_/Y sky130_fd_sc_hd__inv_2
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05829_ _05828_/Q _05852_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_09597_ _09632_/A VGND VGND VPWR VPWR _09597_/Y sky130_fd_sc_hd__inv_2
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08560_/CLK line[112] VGND VGND VPWR VPWR _08548_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[29\] _10867_/Z _10377_/Z _07087_/Z _13597_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[29] sky130_fd_sc_hd__mux4_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11043__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _08478_/Q _08512_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06137__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ _10520_/CLK line[122] VGND VGND VPWR VPWR _10511_/A sky130_fd_sc_hd__dfxtp_1
X_11490_ _11500_/CLK line[58] VGND VGND VPWR VPWR _11490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05041__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11978__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10882__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10441_ _10441_/A _10472_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05976__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[5\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _12570_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08352__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13160_ _13159_/Q _13167_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_10372_ _10384_/CLK line[59] VGND VGND VPWR VPWR _10372_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[8\].TOBUF OVHB\[15\].VALID\[8\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_12111_ _12109_/CLK line[72] VGND VGND VPWR VPWR _12111_/Q sky130_fd_sc_hd__dfxtp_1
X_13091_ _13075_/CLK line[8] VGND VGND VPWR VPWR _13091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12042_ _12042_/A _12047_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[4\].FF OVHB\[3\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[3\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06600__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11218__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12944_ _12943_/Q _12957_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05216__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ _12881_/CLK line[37] VGND VGND VPWR VPWR _12875_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13433__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08527__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11826_ _11825_/Q _11837_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[25\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _09910_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11757_ _11757_/CLK line[38] VGND VGND VPWR VPWR _11757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _10708_/A _10717_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _11687_/Q _11697_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09001__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10792__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13427_ _13439_/CLK line[33] VGND VGND VPWR VPWR _13427_/Q sky130_fd_sc_hd__dfxtp_1
X_10639_ _10627_/CLK line[39] VGND VGND VPWR VPWR _10640_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13358_ _13357_/Q _13377_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12309_ _12311_/CLK line[34] VGND VGND VPWR VPWR _12309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12362__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13289_ _13285_/CLK line[98] VGND VGND VPWR VPWR _13289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12081__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13608__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07850_ _07854_/CLK line[58] VGND VGND VPWR VPWR _07850_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09093__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06801_ _06800_/Q _06832_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_07781_ _07780_/Q _07812_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_04993_ _04992_/Q _05012_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_09520_ _09520_/A _09527_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10032__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06732_ _06740_/CLK line[59] VGND VGND VPWR VPWR _06732_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[7\].TOBUF OVHB\[21\].VALID\[7\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_37_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05126__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[1\].VALID\[6\].FF OVHB\[1\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[1\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10967__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09451_ _09427_/CLK line[8] VGND VGND VPWR VPWR _09451_/Q sky130_fd_sc_hd__dfxtp_1
X_06663_ _06662_/Q _06692_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13343__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05614_ _05632_/CLK line[60] VGND VGND VPWR VPWR _05614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08402_ _08401_/Q _08407_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04965__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09382_ _09381_/Q _09387_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_06594_ _06596_/CLK line[124] VGND VGND VPWR VPWR _06594_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07341__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08333_ _08329_/CLK line[9] VGND VGND VPWR VPWR _08333_/Q sky130_fd_sc_hd__dfxtp_1
X_05545_ _05544_/Q _05572_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12537__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08264_ _08263_/Q _08267_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_05476_ _05476_/CLK line[125] VGND VGND VPWR VPWR _05476_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11798__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12256__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07215_ _07215_/CLK _07216_/X VGND VGND VPWR VPWR _07183_/CLK sky130_fd_sc_hd__dlclkp_1
X_08195_ _08195_/CLK _08196_/X VGND VGND VPWR VPWR _08175_/CLK sky130_fd_sc_hd__dlclkp_1
XDATA\[24\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _09525_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09268__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[29\]_A1 _10377_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07146_ _07111_/A wr VGND VGND VPWR VPWR _07146_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[29\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10207__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07077_ _07111_/A VGND VGND VPWR VPWR _07077_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06028_ _06050_/CLK line[112] VGND VGND VPWR VPWR _06028_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08900__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13518__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12422__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07516__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07979_ _07981_/CLK line[103] VGND VGND VPWR VPWR _07979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09718_ _09717_/Q _09737_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08197__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10990_ _10989_/Q _10997_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09731__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09649_ _09659_/CLK line[98] VGND VGND VPWR VPWR _09650_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13831__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12659_/Q _12677_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11605_/CLK line[99] VGND VGND VPWR VPWR _11611_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12601_/CLK line[35] VGND VGND VPWR VPWR _12591_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _11542_/A _11557_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[13\].TOBUF OVHB\[17\].VALID\[13\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _11479_/CLK line[36] VGND VGND VPWR VPWR _11474_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09178__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13212_ _13211_/Q _13237_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08082__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10424_ _10423_/Q _10437_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13143_ _13163_/CLK line[46] VGND VGND VPWR VPWR _13143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10355_ _10341_/CLK line[37] VGND VGND VPWR VPWR _10355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09906__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13074_ _13074_/A _13097_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_10286_ _10285_/Q _10297_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_12025_ _12019_/CLK line[47] VGND VGND VPWR VPWR _12025_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12332__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[13\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _06270_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09491__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[1\].FF OVHB\[28\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[28\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06330__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13976_ _13979_/A _13979_/B _13979_/C _13979_/D VGND VGND VPWR VPWR _13976_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__09641__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12927_ _12937_/CLK line[75] VGND VGND VPWR VPWR _12927_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[12\].TOBUF OVHB\[10\].VALID\[12\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13163__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08257__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ _12857_/Q _12887_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11809_ _11823_/CLK line[76] VGND VGND VPWR VPWR _11809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12789_ _12803_/CLK line[12] VGND VGND VPWR VPWR _12789_/Q sky130_fd_sc_hd__dfxtp_1
X_05330_ _05332_/CLK line[58] VGND VGND VPWR VPWR _05330_/Q sky130_fd_sc_hd__dfxtp_1
X_05261_ _05260_/Q _05292_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12507__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11411__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07000_ _06999_/Q _07007_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09666__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06505__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05192_ _05214_/CLK line[123] VGND VGND VPWR VPWR _05193_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09816__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08951_ _08947_/CLK line[35] VGND VGND VPWR VPWR _08951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[14\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13338__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07902_ _07902_/A _07917_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13916__A A[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08882_ _08881_/Q _08897_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06240__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07833_ _07837_/CLK line[36] VGND VGND VPWR VPWR _07833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07764_ _07763_/Q _07777_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_04976_ _05152_/A wr VGND VGND VPWR VPWR _04976_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[16\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[12\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _05885_/CLK sky130_fd_sc_hd__clkbuf_4
X_09503_ _09507_/CLK line[46] VGND VGND VPWR VPWR _09503_/Q sky130_fd_sc_hd__dfxtp_1
X_06715_ _06711_/CLK line[37] VGND VGND VPWR VPWR _06715_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10697__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07695_ _07679_/CLK line[101] VGND VGND VPWR VPWR _07695_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13073__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08167__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09434_ _09433_/Q _09457_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06646_ _06645_/Q _06657_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07071__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[3\].FF OVHB\[26\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[26\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _09365_/CLK line[111] VGND VGND VPWR VPWR _09366_/A sky130_fd_sc_hd__dfxtp_1
X_06577_ _06565_/CLK line[102] VGND VGND VPWR VPWR _06577_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11171__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08316_ _08315_/Q _08337_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05528_ _05527_/Q _05537_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_09296_ _09295_/Q _09317_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08247_ _08257_/CLK line[97] VGND VGND VPWR VPWR _08247_/Q sky130_fd_sc_hd__dfxtp_1
X_05459_ _05445_/CLK line[103] VGND VGND VPWR VPWR _05460_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11321__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06415__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08178_ _08177_/Q _08197_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _07117_/CLK line[98] VGND VGND VPWR VPWR _07129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[10\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10140_ _10139_/Q _10157_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08630__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[11\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13248__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[12\].TOBUF OVHB\[30\].VALID\[12\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_10071_ _10073_/CLK line[35] VGND VGND VPWR VPWR _10071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07246__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11346__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13830_ _13830_/CLK _13831_/X VGND VGND VPWR VPWR _13822_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_90_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[4\].TOBUF OVHB\[3\].VALID\[4\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_13761_ _13907_/X wr VGND VGND VPWR VPWR _13761_/X sky130_fd_sc_hd__and2_1
X_10973_ _10977_/CLK line[78] VGND VGND VPWR VPWR _10973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12712_ _12712_/A VGND VGND VPWR VPWR _12712_/Y sky130_fd_sc_hd__inv_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[28\].VALID\[7\].TOBUF OVHB\[28\].VALID\[7\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_13692_ _13907_/X VGND VGND VPWR VPWR _13692_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12643_ _12667_/CLK line[64] VGND VGND VPWR VPWR _12643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13711__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ _12573_/Q _12607_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VOBUF OVHB\[29\].V/Q OVHB\[29\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _11535_/CLK line[74] VGND VGND VPWR VPWR _11525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[5\].FF OVHB\[24\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[24\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11456_ _11455_/Q _11487_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10407_ _10405_/CLK line[75] VGND VGND VPWR VPWR _10407_/Q sky130_fd_sc_hd__dfxtp_1
X_11387_ _11395_/CLK line[11] VGND VGND VPWR VPWR _11387_/Q sky130_fd_sc_hd__dfxtp_1
X_13126_ _13120_/CLK line[24] VGND VGND VPWR VPWR _13127_/A sky130_fd_sc_hd__dfxtp_1
X_10338_ _10337_/Q _10367_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12062__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _13056_/Q _13062_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_10269_ _10277_/CLK line[12] VGND VGND VPWR VPWR _10269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07156__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12008_ _12002_/CLK line[25] VGND VGND VPWR VPWR _12008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12997__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06995__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09371__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[19\]_A0 _10877_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13959_ A_h[5] VGND VGND VPWR VPWR _13964_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06500_ _06499_/Q _06517_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10310__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07480_ _07479_/Q _07497_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05404__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06431_ _06421_/CLK line[35] VGND VGND VPWR VPWR _06431_/Q sky130_fd_sc_hd__dfxtp_1
X_06362_ _06361_/Q _06377_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_09150_ _09149_/Q _09177_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_08101_ _08113_/CLK line[45] VGND VGND VPWR VPWR _08101_/Q sky130_fd_sc_hd__dfxtp_1
X_05313_ _05299_/CLK line[36] VGND VGND VPWR VPWR _05313_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12237__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06293_ _06285_/CLK line[100] VGND VGND VPWR VPWR _06293_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ _09085_/CLK line[109] VGND VGND VPWR VPWR _09081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08032_ _08032_/A _08057_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_05244_ _05243_/Q _05257_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05175_ _05157_/CLK line[101] VGND VGND VPWR VPWR _05175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09546__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09983_ _10011_/CLK line[0] VGND VGND VPWR VPWR _09983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08934_ _08934_/A _08967_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[7\].FF OVHB\[22\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[22\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08865_ _08869_/CLK line[10] VGND VGND VPWR VPWR _08865_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[12\].FF OVHB\[30\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[30\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07816_ _07815_/Q _07847_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12700__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08796_ _08795_/Q _08827_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[12\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07747_ _07773_/CLK line[11] VGND VGND VPWR VPWR _07747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04959_ _04947_/CLK line[2] VGND VGND VPWR VPWR _04960_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07678_ _07677_/Q _07707_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DECH.DEC0.AND1_A_N A_h[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09417_ _09417_/A _09422_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06629_ _06633_/CLK line[12] VGND VGND VPWR VPWR _06629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _09320_/CLK line[89] VGND VGND VPWR VPWR _09348_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VOBUF OVHB\[30\].V/Q OVHB\[30\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XMUX.MUX\[11\] _04948_/Z _05578_/Z _13488_/Z _07118_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[11] sky130_fd_sc_hd__mux4_1
X_09279_ _09278_/Q _09282_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11051__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11310_ _11310_/CLK _11311_/X VGND VGND VPWR VPWR _11302_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06145__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12290_ _12290_/CLK _12291_/X VGND VGND VPWR VPWR _12268_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11986__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11241_ _11311_/A wr VGND VGND VPWR VPWR _11241_/X sky130_fd_sc_hd__and2_1
XOVHB\[1\].VALID\[9\].TOBUF OVHB\[1\].VALID\[9\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[14\].FF OVHB\[20\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[20\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[5\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05984__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08360__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11172_ _11311_/A VGND VGND VPWR VPWR _11172_/Y sky130_fd_sc_hd__inv_2
X_10123_ _10145_/CLK line[64] VGND VGND VPWR VPWR _10123_/Q sky130_fd_sc_hd__dfxtp_1
X_10054_ _10053_/Q _10087_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12610__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13813_ _13812_/Q _13832_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11226__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[20\].VALID\[9\].FF OVHB\[20\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[20\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13744_ _13746_/CLK line[50] VGND VGND VPWR VPWR _13744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10956_ _10930_/CLK line[56] VGND VGND VPWR VPWR _10956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13675_ _13674_/Q _13692_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13441__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10887_ _10886_/Q _10892_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08535__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _12638_/CLK line[51] VGND VGND VPWR VPWR _12626_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12557_ _12556_/Q _12572_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _11500_/CLK line[52] VGND VGND VPWR VPWR _11508_/Q sky130_fd_sc_hd__dfxtp_1
X_12488_ _12490_/CLK line[116] VGND VGND VPWR VPWR _12488_/Q sky130_fd_sc_hd__dfxtp_1
X_11439_ _11439_/A _11452_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05894__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08270__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13109_ _13108_/Q _13132_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_06980_ _06979_/Q _07007_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_05931_ _05929_/CLK line[77] VGND VGND VPWR VPWR _05931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[12\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13616__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08650_ _08650_/CLK _08651_/X VGND VGND VPWR VPWR _08646_/CLK sky130_fd_sc_hd__dlclkp_1
X_05862_ _05861_/Q _05887_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_07601_ _07672_/A wr VGND VGND VPWR VPWR _07601_/X sky130_fd_sc_hd__and2_1
X_08581_ _13921_/X wr VGND VGND VPWR VPWR _08581_/X sky130_fd_sc_hd__and2_1
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05793_ _05799_/CLK line[14] VGND VGND VPWR VPWR _05793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10040__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07532_ _07672_/A VGND VGND VPWR VPWR _07532_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05134__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05712__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10975__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07463_ _07467_/CLK line[0] VGND VGND VPWR VPWR _07463_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13351__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09202_ _09200_/CLK line[22] VGND VGND VPWR VPWR _09202_/Q sky130_fd_sc_hd__dfxtp_1
X_06414_ _06413_/Q _06447_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04973__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05431__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08445__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07394_ _07393_/Q _07427_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_09133_ _09132_/Q _09142_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_06345_ _06353_/CLK line[10] VGND VGND VPWR VPWR _06345_/Q sky130_fd_sc_hd__dfxtp_1
X_06276_ _06275_/Q _06307_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_09064_ _09068_/CLK line[87] VGND VGND VPWR VPWR _09064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05227_ _05253_/CLK line[11] VGND VGND VPWR VPWR _05227_/Q sky130_fd_sc_hd__dfxtp_1
X_08015_ _08014_/Q _08022_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09276__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05158_ _05157_/Q _05187_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13376__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10215__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09966_ _09978_/CLK line[115] VGND VGND VPWR VPWR _09966_/Q sky130_fd_sc_hd__dfxtp_1
X_05089_ _05093_/CLK line[76] VGND VGND VPWR VPWR _05090_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05309__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08917_ _08916_/Q _08932_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09897_ _09897_/A _09912_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13526__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[3\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _12185_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[26\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05606__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08848_ _08850_/CLK line[116] VGND VGND VPWR VPWR _08848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[11\].TOBUF OVHB\[27\].VALID\[11\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07524__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[14\].TOBUF OVHB\[0\].VALID\[14\].FF/Q OVHB\[0\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08779_ _08778_/Q _08792_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_10810_ _10804_/CLK line[117] VGND VGND VPWR VPWR _10810_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].CG clk OVHB\[11\].CGAND/X VGND VGND VPWR VPWR OVHB\[11\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_11790_ _11776_/CLK line[53] VGND VGND VPWR VPWR _11790_/Q sky130_fd_sc_hd__dfxtp_1
X_10741_ _10741_/A _10752_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13460_ _13468_/CLK line[63] VGND VGND VPWR VPWR _13460_/Q sky130_fd_sc_hd__dfxtp_1
X_10672_ _10656_/CLK line[54] VGND VGND VPWR VPWR _10672_/Q sky130_fd_sc_hd__dfxtp_1
X_12411_ _12410_/Q _12432_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_13391_ _13390_/Q _13412_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12342_ _12352_/CLK line[49] VGND VGND VPWR VPWR _12342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _12272_/Q _12292_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09186__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11224_ _11216_/CLK line[50] VGND VGND VPWR VPWR _11224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[10\].TOBUF OVHB\[20\].VALID\[10\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10125__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11155_ _11155_/A _11172_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[25\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10106_ _10100_/CLK line[51] VGND VGND VPWR VPWR _10107_/A sky130_fd_sc_hd__dfxtp_1
X_11086_ _11090_/CLK line[115] VGND VGND VPWR VPWR _11086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12340__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10037_ _10036_/Q _10052_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07434__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[24\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[2\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _11240_/CLK sky130_fd_sc_hd__clkbuf_4
X_11988_ _12002_/CLK line[30] VGND VGND VPWR VPWR _11988_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[16\]_A3 _13589_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13727_ _13907_/X VGND VGND VPWR VPWR _13727_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10939_ _10938_/Q _10962_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13658_ _13682_/CLK line[16] VGND VGND VPWR VPWR _13659_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ _12608_/Q _12642_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_13589_ _13588_/Q _13622_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06130_ _06130_/CLK _06131_/X VGND VGND VPWR VPWR _06108_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_118_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06061_ _13910_/X wr VGND VGND VPWR VPWR _06061_/X sky130_fd_sc_hd__and2_1
XANTENNA__12515__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07609__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05012_ _05152_/A VGND VGND VPWR VPWR _05012_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06513__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09820_ _09834_/CLK line[63] VGND VGND VPWR VPWR _09820_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[9\].TOBUF OVHB\[8\].VALID\[9\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09824__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09751_ _09750_/Q _09772_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06963_ _06962_/Q _06972_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_08702_ _08710_/CLK line[49] VGND VGND VPWR VPWR _08703_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _09140_/CLK sky130_fd_sc_hd__clkbuf_4
X_05914_ _05902_/CLK line[55] VGND VGND VPWR VPWR _05914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09682_ _09694_/CLK line[113] VGND VGND VPWR VPWR _09683_/A sky130_fd_sc_hd__dfxtp_1
X_06894_ _06892_/CLK line[119] VGND VGND VPWR VPWR _06894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08633_ _08632_/Q _08652_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05845_ _05844_/Q _05852_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08564_ _08560_/CLK line[114] VGND VGND VPWR VPWR _08564_/Q sky130_fd_sc_hd__dfxtp_1
X_05776_ _05756_/CLK line[120] VGND VGND VPWR VPWR _05777_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07515_ _07514_/Q _07532_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[6\].CG clk OVHB\[6\].CGAND/X VGND VGND VPWR VPWR OVHB\[6\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13081__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08495_ _08494_/Q _08512_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05799__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08175__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07446_ _07446_/CLK line[115] VGND VGND VPWR VPWR _07447_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[1\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _08055_/CLK sky130_fd_sc_hd__clkbuf_4
X_07377_ _07377_/A _07392_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_09116_ _09116_/CLK line[125] VGND VGND VPWR VPWR _09116_/Q sky130_fd_sc_hd__dfxtp_1
X_06328_ _06320_/CLK line[116] VGND VGND VPWR VPWR _06328_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04932__A1_N A_h[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09047_ _09046_/Q _09072_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_06259_ _06258_/Q _06272_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06423__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05039__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09949_ _09948_/Q _09982_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13256__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12960_ _12962_/CLK line[90] VGND VGND VPWR VPWR _12960_/Q sky130_fd_sc_hd__dfxtp_1
X_11911_ _11910_/Q _11942_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_12891_ _12890_/Q _12922_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_11842_ _11846_/CLK line[91] VGND VGND VPWR VPWR _11842_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[21\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _08755_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[15\].VALID\[4\].TOBUF OVHB\[15\].VALID\[4\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11773_ _11772_/Q _11802_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[24\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11504__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13512_ _13511_/Q _13517_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_10724_ _10728_/CLK line[92] VGND VGND VPWR VPWR _10724_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11801__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13443_ _13439_/CLK line[41] VGND VGND VPWR VPWR _13443_/Q sky130_fd_sc_hd__dfxtp_1
X_10655_ _10654_/Q _10682_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08813__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13374_ _13373_/Q _13377_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10586_ _10594_/CLK line[29] VGND VGND VPWR VPWR _10586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12325_ _12325_/CLK _12326_/X VGND VGND VPWR VPWR _12311_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12256_ _13943_/X wr VGND VGND VPWR VPWR _12256_/X sky130_fd_sc_hd__and2_1
X_11207_ _11311_/A VGND VGND VPWR VPWR _11207_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12187_ _12151_/A VGND VGND VPWR VPWR _12187_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11138_ _11148_/CLK line[16] VGND VGND VPWR VPWR _11138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12070__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11069_ _11068_/Q _11102_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07164__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07742__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05630_ _05632_/CLK line[53] VGND VGND VPWR VPWR _05630_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07461__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05561_ _05560_/Q _05572_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_07300_ _07292_/CLK line[63] VGND VGND VPWR VPWR _07300_/Q sky130_fd_sc_hd__dfxtp_1
X_05492_ _05476_/CLK line[118] VGND VGND VPWR VPWR _05493_/A sky130_fd_sc_hd__dfxtp_1
X_08280_ _08282_/CLK line[127] VGND VGND VPWR VPWR _08280_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05412__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[20\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _08370_/CLK sky130_fd_sc_hd__clkbuf_4
X_07231_ _07230_/Q _07252_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08723__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07162_ _07170_/CLK line[113] VGND VGND VPWR VPWR _07162_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[10\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _05500_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[21\].VALID\[3\].TOBUF OVHB\[21\].VALID\[3\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_06113_ _06112_/Q _06132_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_07093_ _07093_/A _07112_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12245__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07339__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06044_ _06050_/CLK line[114] VGND VGND VPWR VPWR _06044_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07917__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[7\].FF OVHB\[8\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[8\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07636__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09554__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09803_ _09793_/CLK line[41] VGND VGND VPWR VPWR _09804_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07995_ _07994_/Q _08022_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09734_ _09733_/Q _09737_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_06946_ _06960_/CLK line[29] VGND VGND VPWR VPWR _06947_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09665_ _09665_/CLK _09666_/X VGND VGND VPWR VPWR _09659_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[9\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].CGAND_A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06877_ _06877_/A _06902_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13804__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08616_ _13922_/X wr VGND VGND VPWR VPWR _08616_/X sky130_fd_sc_hd__and2_1
XFILLER_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05828_ _05836_/CLK line[30] VGND VGND VPWR VPWR _05828_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09632_/A wr VGND VGND VPWR VPWR _09596_/X sky130_fd_sc_hd__and2_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _13921_/X VGND VGND VPWR VPWR _08547_/Y sky130_fd_sc_hd__inv_2
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05759_ _05758_/Q _05782_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ _08480_/CLK line[80] VGND VGND VPWR VPWR _08478_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[25\].VALID\[14\].FF OVHB\[25\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[25\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07429_ _07428_/Q _07462_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09729__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[6\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10440_ _10466_/CLK line[90] VGND VGND VPWR VPWR _10441_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12155__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10371_ _10370_/Q _10402_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12110_ _12109_/Q _12117_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06153__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13090_ _13089_/Q _13097_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11994__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[9\].TOBUF OVHB\[13\].VALID\[9\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_12041_ _12019_/CLK line[40] VGND VGND VPWR VPWR _12042_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09464__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10403__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12943_ _12937_/CLK line[68] VGND VGND VPWR VPWR _12943_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[9\].FF OVHB\[6\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[6\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12874_ _12873_/Q _12887_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05082__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07712__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ _11823_/CLK line[69] VGND VGND VPWR VPWR _11825_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11234__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06328__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11756_ _11755_/Q _11767_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/CLK line[70] VGND VGND VPWR VPWR _10708_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11691_/CLK line[6] VGND VGND VPWR VPWR _11687_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09639__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13426_ _13425_/Q _13447_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_10638_ _10637_/Q _10647_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08543__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09001__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[22\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13357_ _13347_/CLK line[1] VGND VGND VPWR VPWR _13357_/Q sky130_fd_sc_hd__dfxtp_1
X_10569_ _10571_/CLK line[7] VGND VGND VPWR VPWR _10570_/A sky130_fd_sc_hd__dfxtp_1
X_12308_ _12307_/Q _12327_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06063__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13288_ _13287_/Q _13307_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12239_ _12227_/CLK line[2] VGND VGND VPWR VPWR _12240_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05257__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11409__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06800_ _06802_/CLK line[90] VGND VGND VPWR VPWR _06800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07780_ _07788_/CLK line[26] VGND VGND VPWR VPWR _07780_/Q sky130_fd_sc_hd__dfxtp_1
X_04992_ _05000_/CLK line[17] VGND VGND VPWR VPWR _04992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06731_ _06730_/Q _06762_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09450_ _09450_/A _09457_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08718__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06662_ _06682_/CLK line[27] VGND VGND VPWR VPWR _06662_/Q sky130_fd_sc_hd__dfxtp_1
X_08401_ _08383_/CLK line[40] VGND VGND VPWR VPWR _08401_/Q sky130_fd_sc_hd__dfxtp_1
X_05613_ _05612_/Q _05642_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
X_09381_ _09365_/CLK line[104] VGND VGND VPWR VPWR _09381_/Q sky130_fd_sc_hd__dfxtp_1
X_06593_ _06592_/Q _06622_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11144__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08332_ _08331_/Q _08337_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_05544_ _05568_/CLK line[28] VGND VGND VPWR VPWR _05544_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06238__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05142__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10983__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08263_ _08257_/CLK line[105] VGND VGND VPWR VPWR _08263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05475_ _05474_/Q _05502_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_07214_ _07214_/A _07217_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08453__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08194_ _08194_/A _08197_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_07145_ _07145_/CLK _07146_/X VGND VGND VPWR VPWR _07117_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.MUX\[29\]_A2 _07087_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07069__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06551__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07076_ _07111_/A wr VGND VGND VPWR VPWR _07076_/X sky130_fd_sc_hd__and2_1
X_06027_ _13910_/X VGND VGND VPWR VPWR _06027_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06701__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11319__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10223__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07978_ _07977_/Q _07987_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05317__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09717_ _09721_/CLK line[1] VGND VGND VPWR VPWR _09717_/Q sky130_fd_sc_hd__dfxtp_1
X_06929_ _06923_/CLK line[7] VGND VGND VPWR VPWR _06929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13534__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09648_ _09648_/A _09667_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08628__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[13\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[13\].VALID\[14\].TOBUF OVHB\[13\].VALID\[14\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[1\].FF OVHB\[15\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[15\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13831__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09577_/CLK line[66] VGND VGND VPWR VPWR _09580_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11609_/Q _11627_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12589_/Q _12607_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06726__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05052__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[10\].FF OVHB\[31\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[31\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10893__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11535_/CLK line[67] VGND VGND VPWR VPWR _11542_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[17\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ _11471_/Q _11487_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ _13213_/CLK line[77] VGND VGND VPWR VPWR _13211_/Q sky130_fd_sc_hd__dfxtp_1
X_10423_ _10405_/CLK line[68] VGND VGND VPWR VPWR _10423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[0\].TOBUF OVHB\[3\].VALID\[0\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13142_ _13141_/Q _13167_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_10354_ _10353_/Q _10367_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[28\].VALID\[3\].TOBUF OVHB\[28\].VALID\[3\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13709__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13073_ _13075_/CLK line[14] VGND VGND VPWR VPWR _13074_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10285_ _10277_/CLK line[5] VGND VGND VPWR VPWR _10285_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09194__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ _12023_/Q _12047_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09772__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10133__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09491__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VOBUF OVHB\[25\].V/Q OVHB\[25\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_93_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05227__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13975_ _13979_/C _13979_/B _13979_/A _13979_/D VGND VGND VPWR VPWR _13975_/X sky130_fd_sc_hd__and4b_4
XOVHB\[21\].VALID\[12\].FF OVHB\[21\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[21\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12926_ _12925_/Q _12957_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07442__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12857_ _12881_/CLK line[43] VGND VGND VPWR VPWR _12857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[8\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06058__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11808_ _11807_/Q _11837_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_12788_ _12788_/A _12817_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11899__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11739_ _11757_/CLK line[44] VGND VGND VPWR VPWR _11739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09369__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09947__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05260_ _05278_/CLK line[26] VGND VGND VPWR VPWR _05260_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[3\].FF OVHB\[13\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[13\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05191_ _05191_/A _05222_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_13409_ _13409_/A _13412_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10308__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[7\].FF OVHB\[30\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[30\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09666__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08950_ _08949_/Q _08967_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12523__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[14\].FF OVHB\[11\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[11\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07617__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07901_ _07905_/CLK line[67] VGND VGND VPWR VPWR _07902_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[20\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08881_ _08869_/CLK line[3] VGND VGND VPWR VPWR _08881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07832_ _07832_/A _07847_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09832__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07763_ _07773_/CLK line[4] VGND VGND VPWR VPWR _07763_/Q sky130_fd_sc_hd__dfxtp_1
X_04975_ _04975_/CLK _04976_/X VGND VGND VPWR VPWR _04947_/CLK sky130_fd_sc_hd__dlclkp_1
X_09502_ _09502_/A _09527_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_06714_ _06713_/Q _06727_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07694_ _07694_/A _07707_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09433_ _09427_/CLK line[14] VGND VGND VPWR VPWR _09433_/Q sky130_fd_sc_hd__dfxtp_1
X_06645_ _06633_/CLK line[5] VGND VGND VPWR VPWR _06645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11452__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09364_ _09364_/A _09387_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_06576_ _06575_/Q _06587_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_08315_ _08329_/CLK line[15] VGND VGND VPWR VPWR _08315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11171__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05527_ _05519_/CLK line[6] VGND VGND VPWR VPWR _05527_/Q sky130_fd_sc_hd__dfxtp_1
X_09295_ _09307_/CLK line[79] VGND VGND VPWR VPWR _09295_/Q sky130_fd_sc_hd__dfxtp_1
X_08246_ _08245_/Q _08267_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08183__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05458_ _05457_/Q _05467_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[8\].FF OVHB\[29\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[29\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08177_ _08175_/CLK line[65] VGND VGND VPWR VPWR _08177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05389_ _05391_/CLK line[71] VGND VGND VPWR VPWR _05389_/Q sky130_fd_sc_hd__dfxtp_1
X_07128_ _07127_/Q _07147_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12433__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07059_ _07043_/CLK line[66] VGND VGND VPWR VPWR _07060_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[11\].VALID\[5\].FF OVHB\[11\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[11\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06431__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10070_ _10069_/Q _10087_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11049__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11627__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09742__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11346__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10888__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13264__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13760_ _13760_/CLK _13761_/X VGND VGND VPWR VPWR _13746_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08358__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10972_ _10971_/Q _10997_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].VALID\[5\].TOBUF OVHB\[1\].VALID\[5\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_12711_ _12712_/A wr VGND VGND VPWR VPWR _12711_/X sky130_fd_sc_hd__and2_1
X_13691_ _13907_/X wr VGND VGND VPWR VPWR _13691_/X sky130_fd_sc_hd__and2_1
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ _12712_/A VGND VGND VPWR VPWR _12642_/Y sky130_fd_sc_hd__inv_2
XOVHB\[26\].VALID\[8\].TOBUF OVHB\[26\].VALID\[8\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_31_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12608__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12573_ _12601_/CLK line[32] VGND VGND VPWR VPWR _12573_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11512__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08093__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _11523_/Q _11557_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06606__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11455_ _11479_/CLK line[42] VGND VGND VPWR VPWR _11455_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07287__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10406_ _10405_/Q _10437_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08821__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11386_ _11385_/Q _11417_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13439__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13125_ _13125_/A _13132_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_10337_ _10341_/CLK line[43] VGND VGND VPWR VPWR _10337_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[19\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12921__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13056_ _13050_/CLK line[120] VGND VGND VPWR VPWR _13056_/Q sky130_fd_sc_hd__dfxtp_1
X_10268_ _10267_/Q _10297_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12007_ _12006_/Q _12012_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10199_ _10217_/CLK line[108] VGND VGND VPWR VPWR _10199_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10798__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13174__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08268__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[19\]_A1 _10387_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13958_ A_h[4] VGND VGND VPWR VPWR _13958_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07172__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12909_ _12908_/Q _12922_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_13889_ _13888_/Q _13902_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[30\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _11625_/CLK sky130_fd_sc_hd__clkbuf_4
X_06430_ _06429_/Q _06447_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06361_ _06353_/CLK line[3] VGND VGND VPWR VPWR _06361_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11422__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09099__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08100_ _08100_/A _08127_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_05312_ _05312_/A _05327_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09080_ _09080_/A _09107_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_06292_ _06292_/A _06307_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08581__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05420__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08031_ _08033_/CLK line[13] VGND VGND VPWR VPWR _08032_/A sky130_fd_sc_hd__dfxtp_1
X_05243_ _05253_/CLK line[4] VGND VGND VPWR VPWR _05243_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10038__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08731__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05174_ _05173_/Q _05187_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13349__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12253__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13927__A A[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09982_ _09912_/A VGND VGND VPWR VPWR _09982_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07347__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08933_ _08947_/CLK line[32] VGND VGND VPWR VPWR _08934_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[11\].TOBUF OVHB\[7\].VALID\[11\].FF/Q OVHB\[7\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_08864_ _08863_/Q _08897_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07815_ _07837_/CLK line[42] VGND VGND VPWR VPWR _07815_/Q sky130_fd_sc_hd__dfxtp_1
X_08795_ _08823_/CLK line[106] VGND VGND VPWR VPWR _08795_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10501__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07746_ _07745_/Q _07777_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_04958_ _04957_/Q _04977_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07082__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08756__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07677_ _07679_/CLK line[107] VGND VGND VPWR VPWR _07677_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13812__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09416_ _09414_/CLK line[120] VGND VGND VPWR VPWR _09417_/A sky130_fd_sc_hd__dfxtp_1
X_06628_ _06627_/Q _06657_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08906__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09347_ _09346_/Q _09352_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_06559_ _06565_/CLK line[108] VGND VGND VPWR VPWR _06560_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12428__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09278_ _09256_/CLK line[57] VGND VGND VPWR VPWR _09278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05330__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08229_ _08228_/Q _08232_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[10\].TOBUF OVHB\[0\].VALID\[10\].FF/Q OVHB\[0\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_11240_ _11240_/CLK _11241_/X VGND VGND VPWR VPWR _11216_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12163__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11171_ _11311_/A wr VGND VGND VPWR VPWR _11171_/X sky130_fd_sc_hd__and2_1
XFILLER_136_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07257__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10122_ _10192_/A VGND VGND VPWR VPWR _10122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06161__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10053_ _10073_/CLK line[32] VGND VGND VPWR VPWR _10053_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10261__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09472__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10411__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08088__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13812_ _13822_/CLK line[81] VGND VGND VPWR VPWR _13812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05505__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13743_ _13742_/Q _13762_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_10955_ _10954_/Q _10962_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13674_ _13682_/CLK line[18] VGND VGND VPWR VPWR _13674_/Q sky130_fd_sc_hd__dfxtp_1
X_10886_ _10872_/CLK line[24] VGND VGND VPWR VPWR _10886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07720__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12338__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12625_ _12624_/Q _12642_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06336__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12556_ _12560_/CLK line[19] VGND VGND VPWR VPWR _12556_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _11506_/Q _11522_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12487_/A _12502_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10436__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09647__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11438_ _11440_/CLK line[20] VGND VGND VPWR VPWR _11439_/A sky130_fd_sc_hd__dfxtp_1
X_11369_ _11368_/Q _11382_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06071__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13108_ _13120_/CLK line[30] VGND VGND VPWR VPWR _13108_/Q sky130_fd_sc_hd__dfxtp_1
X_05930_ _05929_/Q _05957_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12801__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _13038_/Q _13062_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05861_ _05871_/CLK line[45] VGND VGND VPWR VPWR _05861_/Q sky130_fd_sc_hd__dfxtp_1
X_07600_ _07600_/CLK _07601_/X VGND VGND VPWR VPWR _07572_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13482__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08580_ _08580_/CLK _08581_/X VGND VGND VPWR VPWR _08560_/CLK sky130_fd_sc_hd__dlclkp_1
X_05792_ _05791_/Q _05817_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_07531_ _07672_/A wr VGND VGND VPWR VPWR _07531_/X sky130_fd_sc_hd__and2_1
XOVHB\[2\].VALID\[0\].FF OVHB\[2\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[2\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[13\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07462_ _13918_/X VGND VGND VPWR VPWR _07462_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06096__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09201_ _09200_/Q _09212_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[5\].TOBUF OVHB\[8\].VALID\[5\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_06413_ _06421_/CLK line[32] VGND VGND VPWR VPWR _06413_/Q sky130_fd_sc_hd__dfxtp_1
X_07393_ _07393_/CLK line[96] VGND VGND VPWR VPWR _07393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11152__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09132_ _09116_/CLK line[118] VGND VGND VPWR VPWR _09132_/Q sky130_fd_sc_hd__dfxtp_1
X_06344_ _06343_/Q _06377_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06246__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10991__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09063_ _09063_/A _09072_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_06275_ _06285_/CLK line[106] VGND VGND VPWR VPWR _06275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08014_ _08000_/CLK line[119] VGND VGND VPWR VPWR _08014_/Q sky130_fd_sc_hd__dfxtp_1
X_05226_ _05225_/Q _05257_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08461__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[14\].FF OVHB\[2\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[2\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13079__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13657__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05157_ _05157_/CLK line[107] VGND VGND VPWR VPWR _05157_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[12\].TOBUF OVHB\[23\].VALID\[12\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13376__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09965_ _09965_/A _09982_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_05088_ _05087_/Q _05117_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_08916_ _08922_/CLK line[19] VGND VGND VPWR VPWR _08916_/Q sky130_fd_sc_hd__dfxtp_1
X_09896_ _09908_/CLK line[83] VGND VGND VPWR VPWR _09897_/A sky130_fd_sc_hd__dfxtp_1
X_08847_ _08846_/Q _08862_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11327__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08778_ _08762_/CLK line[84] VGND VGND VPWR VPWR _08778_/Q sky130_fd_sc_hd__dfxtp_1
X_07729_ _07728_/Q _07742_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13542__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10740_ _10728_/CLK line[85] VGND VGND VPWR VPWR _10741_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08636__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10671_ _10670_/Q _10682_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12410_ _12414_/CLK line[95] VGND VGND VPWR VPWR _12410_/Q sky130_fd_sc_hd__dfxtp_1
X_13390_ _13394_/CLK line[31] VGND VGND VPWR VPWR _13390_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05060__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[2\].FF OVHB\[0\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[0\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12341_ _12340_/Q _12362_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05995__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12272_ _12268_/CLK line[17] VGND VGND VPWR VPWR _12272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[15\].VALID\[0\].TOBUF OVHB\[15\].VALID\[0\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_11223_ _11222_/Q _11242_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ _11148_/CLK line[18] VGND VGND VPWR VPWR _11155_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[12\].FF OVHB\[26\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[26\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13717__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10105_ _10105_/A _10122_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11085_ _11084_/Q _11102_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10036_ _10042_/CLK line[19] VGND VGND VPWR VPWR _10036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10141__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05235__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[24\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13452__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ _11986_/Q _12012_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_13726_ _13907_/X wr VGND VGND VPWR VPWR _13726_/X sky130_fd_sc_hd__and2_1
X_10938_ _10930_/CLK line[62] VGND VGND VPWR VPWR _10938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07450__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12068__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13657_ _13907_/X VGND VGND VPWR VPWR _13657_/Y sky130_fd_sc_hd__inv_2
X_10869_ _10868_/Q _10892_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ _12638_/CLK line[48] VGND VGND VPWR VPWR _12608_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13588_ _13598_/CLK line[112] VGND VGND VPWR VPWR _13588_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[14\].FF OVHB\[16\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[16\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12539_ _12538_/Q _12572_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11700__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09377__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06060_ _06060_/CLK _06061_/X VGND VGND VPWR VPWR _06050_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_67_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05011_ _05152_/A wr VGND VGND VPWR VPWR _05011_/X sky130_fd_sc_hd__and2_1
XANTENNA__10316__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13627__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12531__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06962_ _06960_/CLK line[22] VGND VGND VPWR VPWR _06962_/Q sky130_fd_sc_hd__dfxtp_1
X_09750_ _09760_/CLK line[31] VGND VGND VPWR VPWR _09750_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07625__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08701_ _08700_/Q _08722_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_05913_ _05912_/Q _05922_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_09681_ _09680_/Q _09702_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_06893_ _06892_/Q _06902_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08632_ _08646_/CLK line[17] VGND VGND VPWR VPWR _08632_/Q sky130_fd_sc_hd__dfxtp_1
X_05844_ _05836_/CLK line[23] VGND VGND VPWR VPWR _05844_/Q sky130_fd_sc_hd__dfxtp_1
X_08563_ _08562_/Q _08582_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_05775_ _05774_/Q _05782_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07514_ _07518_/CLK line[18] VGND VGND VPWR VPWR _07514_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04984__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08494_ _08480_/CLK line[82] VGND VGND VPWR VPWR _08494_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07360__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07445_ _07444_/Q _07462_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ _07380_/CLK line[83] VGND VGND VPWR VPWR _07377_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09115_ _09114_/Q _09142_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[11\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06327_ _06327_/A _06342_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12706__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09287__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08191__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09046_ _09068_/CLK line[93] VGND VGND VPWR VPWR _09046_/Q sky130_fd_sc_hd__dfxtp_1
X_06258_ _06244_/CLK line[84] VGND VGND VPWR VPWR _06258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05209_ _05209_/A _05222_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_06189_ _06188_/Q _06202_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12291__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[0\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12441__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09948_ _09978_/CLK line[112] VGND VGND VPWR VPWR _09948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07535__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11057__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09879_ _09878_/Q _09912_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11910_ _11934_/CLK line[122] VGND VGND VPWR VPWR _11910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12890_ _12902_/CLK line[58] VGND VGND VPWR VPWR _12890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09750__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ _11840_/Q _11872_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11772_ _11776_/CLK line[59] VGND VGND VPWR VPWR _11772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08366__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[5\].TOBUF OVHB\[13\].VALID\[5\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_41_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[30\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13511_ _13497_/CLK line[72] VGND VGND VPWR VPWR _13511_/Q sky130_fd_sc_hd__dfxtp_1
X_10723_ _10722_/Q _10752_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12466__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10654_ _10656_/CLK line[60] VGND VGND VPWR VPWR _10654_/Q sky130_fd_sc_hd__dfxtp_1
X_13442_ _13441_/Q _13447_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12616__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13373_ _13347_/CLK line[9] VGND VGND VPWR VPWR _13373_/Q sky130_fd_sc_hd__dfxtp_1
X_10585_ _10584_/Q _10612_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12324_ _12324_/A _12327_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06614__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12255_ _12255_/CLK _12256_/X VGND VGND VPWR VPWR _12227_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09925__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11206_ _11311_/A wr VGND VGND VPWR VPWR _11206_/X sky130_fd_sc_hd__and2_1
X_12186_ _12151_/A wr VGND VGND VPWR VPWR _12186_/X sky130_fd_sc_hd__and2_1
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11137_ _11311_/A VGND VGND VPWR VPWR _11137_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11068_ _11090_/CLK line[112] VGND VGND VPWR VPWR _11068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ _10018_/Q _10052_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13182__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08276__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05560_ _05568_/CLK line[21] VGND VGND VPWR VPWR _05560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13709_ _13701_/CLK line[34] VGND VGND VPWR VPWR _13709_/Q sky130_fd_sc_hd__dfxtp_1
X_05491_ _05490_/Q _05502_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_07230_ _07232_/CLK line[31] VGND VGND VPWR VPWR _07230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07161_ _07160_/Q _07182_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[10\].FF OVHB\[22\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[22\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11430__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06112_ _06108_/CLK line[17] VGND VGND VPWR VPWR _06112_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06524__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07092_ _07098_/CLK line[81] VGND VGND VPWR VPWR _07093_/A sky130_fd_sc_hd__dfxtp_1
X_06043_ _06042_/Q _06062_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10046__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13357__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09802_ _09801_/Q _09807_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07994_ _08000_/CLK line[124] VGND VGND VPWR VPWR _07994_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[1\].FF OVHB\[23\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[23\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09733_ _09721_/CLK line[9] VGND VGND VPWR VPWR _09733_/Q sky130_fd_sc_hd__dfxtp_1
X_06945_ _06944_/Q _06972_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09664_ _09664_/A _09667_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06876_ _06892_/CLK line[125] VGND VGND VPWR VPWR _06877_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[28\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08615_ _08615_/CLK _08616_/X VGND VGND VPWR VPWR _08609_/CLK sky130_fd_sc_hd__dlclkp_1
X_05827_ _05827_/A _05852_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_09595_ _09595_/CLK _09596_/X VGND VGND VPWR VPWR _09577_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11605__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[29\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[12\].FF OVHB\[12\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[12\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _13921_/X wr VGND VGND VPWR VPWR _08546_/X sky130_fd_sc_hd__and2_1
X_05758_ _05756_/CLK line[126] VGND VGND VPWR VPWR _05758_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07090__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05603__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ _13921_/X VGND VGND VPWR VPWR _08477_/Y sky130_fd_sc_hd__inv_2
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05689_ _05688_/Q _05712_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13820__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ _07446_/CLK line[112] VGND VGND VPWR VPWR _07428_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08914__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[3\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07359_ _07358_/Q _07392_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[6\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10370_ _10384_/CLK line[58] VGND VGND VPWR VPWR _10370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[13\].VALID\[10\].TOBUF OVHB\[13\].VALID\[10\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_09029_ _09005_/CLK line[71] VGND VGND VPWR VPWR _09030_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[14\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12040_ _12039_/Q _12047_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12171__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07265__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ _12941_/Q _12957_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09480__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12873_ _12881_/CLK line[36] VGND VGND VPWR VPWR _12873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[21\].VALID\[3\].FF OVHB\[21\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[21\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11824_ _11823_/Q _11837_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05513__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11755_ _11757_/CLK line[37] VGND VGND VPWR VPWR _11755_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13730__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10705_/Q _10717_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11686_ _11685_/Q _11697_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[21\].VOBUF OVHB\[21\].V/Q OVHB\[21\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__12346__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13425_ _13439_/CLK line[47] VGND VGND VPWR VPWR _13425_/Q sky130_fd_sc_hd__dfxtp_1
X_10637_ _10627_/CLK line[38] VGND VGND VPWR VPWR _10637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[24\].CG clk OVHB\[24\].CGAND/X VGND VGND VPWR VPWR OVHB\[24\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10568_ _10568_/A _10577_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_13356_ _13355_/Q _13377_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12307_ _12311_/CLK line[33] VGND VGND VPWR VPWR _12307_/Q sky130_fd_sc_hd__dfxtp_1
X_13287_ _13285_/CLK line[97] VGND VGND VPWR VPWR _13287_/Q sky130_fd_sc_hd__dfxtp_1
X_10499_ _10473_/CLK line[103] VGND VGND VPWR VPWR _10499_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09655__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12238_ _12237_/Q _12257_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12169_ _12177_/CLK line[98] VGND VGND VPWR VPWR _12169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[7\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04991_ _04990_/Q _05012_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_06730_ _06740_/CLK line[58] VGND VGND VPWR VPWR _06730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09390__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07903__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06661_ _06660_/Q _06692_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05612_ _05632_/CLK line[59] VGND VGND VPWR VPWR _05612_/Q sky130_fd_sc_hd__dfxtp_1
X_08400_ _08399_/Q _08407_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_09380_ _09379_/Q _09387_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06592_ _06596_/CLK line[123] VGND VGND VPWR VPWR _06592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08331_ _08329_/CLK line[8] VGND VGND VPWR VPWR _08331_/Q sky130_fd_sc_hd__dfxtp_1
X_05543_ _05542_/Q _05572_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[14\].FF OVHB\[7\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[7\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08262_ _08261_/Q _08267_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_05474_ _05476_/CLK line[124] VGND VGND VPWR VPWR _05474_/Q sky130_fd_sc_hd__dfxtp_1
X_07213_ _07183_/CLK line[9] VGND VGND VPWR VPWR _07214_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08193_ _08175_/CLK line[73] VGND VGND VPWR VPWR _08194_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11160__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07144_ _07143_/Q _07147_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06254__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[29\]_A3 _13597_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06832__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07075_ _07075_/CLK _07076_/X VGND VGND VPWR VPWR _07043_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[9\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06551__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09565__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06026_ _13910_/X wr VGND VGND VPWR VPWR _06026_/X sky130_fd_sc_hd__and2_1
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13087__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07977_ _07981_/CLK line[102] VGND VGND VPWR VPWR _07977_/Q sky130_fd_sc_hd__dfxtp_1
X_09716_ _09715_/Q _09737_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_06928_ _06927_/Q _06937_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07813__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09647_ _09659_/CLK line[97] VGND VGND VPWR VPWR _09648_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06859_ _06839_/CLK line[103] VGND VGND VPWR VPWR _06860_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11335__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06429__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09578_ _09578_/A _09597_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08541_/CLK line[98] VGND VGND VPWR VPWR _08530_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06726__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _11540_/A _11557_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[18\].VALID\[6\].FF OVHB\[18\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[18\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ _11479_/CLK line[35] VGND VGND VPWR VPWR _11471_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11070__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13209_/Q _13237_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_10422_ _10421_/Q _10437_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10353_ _10341_/CLK line[36] VGND VGND VPWR VPWR _10353_/Q sky130_fd_sc_hd__dfxtp_1
X_13141_ _13163_/CLK line[45] VGND VGND VPWR VPWR _13141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[1\].VALID\[1\].TOBUF OVHB\[1\].VALID\[1\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_136_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13072_ _13071_/Q _13097_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_10284_ _10283_/Q _10297_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[4\].TOBUF OVHB\[26\].VALID\[4\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_12023_ _12019_/CLK line[46] VGND VGND VPWR VPWR _12023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08819__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13974_ _13979_/C _13979_/A _13979_/B _13979_/D VGND VGND VPWR VPWR _13974_/X sky130_fd_sc_hd__and4bb_4
X_12925_ _12937_/CLK line[74] VGND VGND VPWR VPWR _12925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11245__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12856_ _12855_/Q _12887_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].CGAND_A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05243__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11807_ _11823_/CLK line[75] VGND VGND VPWR VPWR _11807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13460__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12787_ _12803_/CLK line[11] VGND VGND VPWR VPWR _12788_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08554__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11738_ _11737_/Q _11767_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].CGAND _13932_/X wr VGND VGND VPWR VPWR OVHB\[28\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__12076__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11669_ _11691_/CLK line[12] VGND VGND VPWR VPWR _11669_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13394_/CLK line[25] VGND VGND VPWR VPWR _13409_/A sky130_fd_sc_hd__dfxtp_1
X_05190_ _05214_/CLK line[122] VGND VGND VPWR VPWR _05191_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[0\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].V OVHB\[2\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[2\].V/Q sky130_fd_sc_hd__dfrtp_1
X_13339_ _13339_/A _13342_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[16\].VALID\[8\].FF OVHB\[16\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[16\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06802__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07900_ _07900_/A _07917_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10324__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08880_ _08879_/Q _08897_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05418__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07831_ _07837_/CLK line[35] VGND VGND VPWR VPWR _07832_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13635__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08729__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07762_ _07761_/Q _07777_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_04974_ _04973_/Q _04977_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07633__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09501_ _09507_/CLK line[45] VGND VGND VPWR VPWR _09502_/A sky130_fd_sc_hd__dfxtp_1
X_06713_ _06711_/CLK line[36] VGND VGND VPWR VPWR _06713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07693_ _07679_/CLK line[100] VGND VGND VPWR VPWR _07694_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06644_ _06643_/Q _06657_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_09432_ _09431_/Q _09457_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05153__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09363_ _09365_/CLK line[110] VGND VGND VPWR VPWR _09364_/A sky130_fd_sc_hd__dfxtp_1
X_06575_ _06565_/CLK line[101] VGND VGND VPWR VPWR _06575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ _08313_/Q _08337_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_05526_ _05525_/Q _05537_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04992__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09294_ _09293_/Q _09317_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_08245_ _08257_/CLK line[111] VGND VGND VPWR VPWR _08245_/Q sky130_fd_sc_hd__dfxtp_1
X_05457_ _05445_/CLK line[102] VGND VGND VPWR VPWR _05457_/Q sky130_fd_sc_hd__dfxtp_1
X_08176_ _08176_/A _08197_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_05388_ _05387_/Q _05397_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
X_07127_ _07117_/CLK line[97] VGND VGND VPWR VPWR _07127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09295__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07808__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07058_ _07057_/Q _07077_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06009_ _06023_/CLK line[98] VGND VGND VPWR VPWR _06009_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10234__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05328__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[3\].VALID\[12\].FF OVHB\[3\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[3\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07543__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10971_ _10977_/CLK line[77] VGND VGND VPWR VPWR _10971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _12710_/CLK _12711_/X VGND VGND VPWR VPWR _12708_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06159__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13690_ _13690_/CLK _13691_/X VGND VGND VPWR VPWR _13682_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05641__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _12712_/A wr VGND VGND VPWR VPWR _12641_/X sky130_fd_sc_hd__and2_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[9\].TOBUF OVHB\[24\].VALID\[9\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _12712_/A VGND VGND VPWR VPWR _12572_/Y sky130_fd_sc_hd__inv_2
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10409__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11523_ _11535_/CLK line[64] VGND VGND VPWR VPWR _11523_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11454_ _11453_/Q _11487_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12624__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10405_ _10405_/CLK line[74] VGND VGND VPWR VPWR _10405_/Q sky130_fd_sc_hd__dfxtp_1
X_11385_ _11395_/CLK line[10] VGND VGND VPWR VPWR _11385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07718__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[9\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _13655_/CLK sky130_fd_sc_hd__clkbuf_4
X_13124_ _13120_/CLK line[23] VGND VGND VPWR VPWR _13125_/A sky130_fd_sc_hd__dfxtp_1
X_10336_ _10335_/Q _10367_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12921__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10267_ _10277_/CLK line[11] VGND VGND VPWR VPWR _10267_/Q sky130_fd_sc_hd__dfxtp_1
X_13055_ _13054_/Q _13062_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09933__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05816__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12006_ _12002_/CLK line[24] VGND VGND VPWR VPWR _12006_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ _10197_/Q _10227_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[21\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13957_ _13950_/A _13950_/B _13950_/C _13957_/D VGND VGND VPWR VPWR _13957_/X sky130_fd_sc_hd__and4_4
XANTENNA_MUX.MUX\[19\]_A2 _07097_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12908_ _12902_/CLK line[52] VGND VGND VPWR VPWR _12908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06069__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13888_ _13882_/CLK line[116] VGND VGND VPWR VPWR _13888_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[10\].FF OVHB\[27\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[27\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12839_ _12839_/A _12852_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13190__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06360_ _06359_/Q _06377_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08284__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08862__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05311_ _05299_/CLK line[35] VGND VGND VPWR VPWR _05312_/A sky130_fd_sc_hd__dfxtp_1
X_06291_ _06285_/CLK line[99] VGND VGND VPWR VPWR _06292_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[29\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _10995_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_30_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08581__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08030_ _08030_/A _08057_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_05242_ _05242_/A _05257_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[12\].TOBUF OVHB\[3\].VALID\[12\].FF/Q OVHB\[3\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_128_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05173_ _05157_/CLK line[100] VGND VGND VPWR VPWR _05173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06532__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[8\].TOBUF OVHB\[30\].VALID\[8\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_09981_ _09912_/A wr VGND VGND VPWR VPWR _09981_/X sky130_fd_sc_hd__and2_1
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08932_ _13923_/X VGND VGND VPWR VPWR _08932_/Y sky130_fd_sc_hd__inv_2
XOVHB\[9\].VALID\[1\].FF OVHB\[9\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[9\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[1\].TOBUF OVHB\[8\].VALID\[1\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05148__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09843__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10989__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08863_ _08869_/CLK line[0] VGND VGND VPWR VPWR _08863_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[12\].FF OVHB\[17\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[17\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13365__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07814_ _07813_/Q _07847_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08459__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08794_ _08793_/Q _08827_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07745_ _07773_/CLK line[10] VGND VGND VPWR VPWR _07745_/Q sky130_fd_sc_hd__dfxtp_1
X_04957_ _04947_/CLK line[1] VGND VGND VPWR VPWR _04957_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08756__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07676_ _07675_/Q _07707_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[14\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09415_ _09414_/Q _09422_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_06627_ _06633_/CLK line[11] VGND VGND VPWR VPWR _06627_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11613__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[1\]_A0 _04958_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06707__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06558_ _06558_/A _06587_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_09346_ _09320_/CLK line[88] VGND VGND VPWR VPWR _09346_/Q sky130_fd_sc_hd__dfxtp_1
X_05509_ _05519_/CLK line[12] VGND VGND VPWR VPWR _05509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09277_ _09277_/A _09282_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_06489_ _06489_/CLK line[76] VGND VGND VPWR VPWR _06489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08922__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08228_ _08208_/CLK line[89] VGND VGND VPWR VPWR _08228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[27\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08159_ _08158_/Q _08162_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[28\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _10610_/CLK sky130_fd_sc_hd__clkbuf_4
X_11170_ _11170_/CLK _11171_/X VGND VGND VPWR VPWR _11148_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_101_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[24\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10121_ _10192_/A wr VGND VGND VPWR VPWR _10121_/X sky130_fd_sc_hd__and2_1
XFILLER_136_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[18\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _07740_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10542__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05058__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10052_ _10192_/A VGND VGND VPWR VPWR _10052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10899__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10261__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13275__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07273__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13811_ _13810_/Q _13832_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[7\].VALID\[3\].FF OVHB\[7\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[7\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13742_ _13746_/CLK line[49] VGND VGND VPWR VPWR _13742_/Q sky130_fd_sc_hd__dfxtp_1
X_10954_ _10930_/CLK line[55] VGND VGND VPWR VPWR _10954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13673_ _13672_/Q _13692_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11523__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10885_ _10885_/A _10892_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12624_ _12638_/CLK line[50] VGND VGND VPWR VPWR _12624_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05521__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _12554_/Q _12572_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10717__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _11500_/CLK line[51] VGND VGND VPWR VPWR _11506_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08832__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12490_/CLK line[115] VGND VGND VPWR VPWR _12487_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10436__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12354__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11437_ _11436_/Q _11452_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07448__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11368_ _11370_/CLK line[116] VGND VGND VPWR VPWR _11368_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[14\].TOBUF OVHB\[26\].VALID\[14\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_13107_ _13106_/Q _13132_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_10319_ _10319_/A _10332_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09663__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11299_ _11298_/Q _11312_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_13038_ _13050_/CLK line[126] VGND VGND VPWR VPWR _13038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05860_ _05860_/A _05887_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10602__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07183__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _07355_/CLK sky130_fd_sc_hd__clkbuf_4
X_05791_ _05799_/CLK line[13] VGND VGND VPWR VPWR _05791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ _07530_/CLK _07531_/X VGND VGND VPWR VPWR _07518_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06377__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07911__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07461_ _13918_/X wr VGND VGND VPWR VPWR _07461_/X sky130_fd_sc_hd__and2_1
XANTENNA__12529__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06096__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06412_ _06551_/A VGND VGND VPWR VPWR _06412_/Y sky130_fd_sc_hd__inv_2
X_09200_ _09200_/CLK line[21] VGND VGND VPWR VPWR _09200_/Q sky130_fd_sc_hd__dfxtp_1
X_07392_ _13918_/X VGND VGND VPWR VPWR _07392_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[6\].VALID\[6\].TOBUF OVHB\[6\].VALID\[6\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[5\].FF OVHB\[5\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[5\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09131_ _09131_/A _09142_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_06343_ _06353_/CLK line[0] VGND VGND VPWR VPWR _06343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09838__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09062_ _09068_/CLK line[86] VGND VGND VPWR VPWR _09063_/A sky130_fd_sc_hd__dfxtp_1
X_06274_ _06273_/Q _06307_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_05225_ _05253_/CLK line[10] VGND VGND VPWR VPWR _05225_/Q sky130_fd_sc_hd__dfxtp_1
X_08013_ _08012_/Q _08022_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12264__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13938__A A[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07358__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06262__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05156_ _05155_/Q _05187_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[29\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09964_ _09978_/CLK line[114] VGND VGND VPWR VPWR _09965_/A sky130_fd_sc_hd__dfxtp_1
X_05087_ _05093_/CLK line[75] VGND VGND VPWR VPWR _05087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09573__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08915_ _08914_/Q _08932_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
X_09895_ _09894_/Q _09912_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10512__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08189__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08846_ _08850_/CLK line[115] VGND VGND VPWR VPWR _08846_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07671__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08777_ _08776_/Q _08792_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_05989_ _05988_/Q _05992_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07728_ _07724_/CLK line[116] VGND VGND VPWR VPWR _07728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07821__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12439__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _06970_/CLK sky130_fd_sc_hd__clkbuf_4
X_07659_ _07658_/Q _07672_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11343__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06437__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10670_ _10656_/CLK line[53] VGND VGND VPWR VPWR _10670_/Q sky130_fd_sc_hd__dfxtp_1
X_09329_ _09328_/Q _09352_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09748__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12340_ _12352_/CLK line[63] VGND VGND VPWR VPWR _12340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12271_ _12270_/Q _12292_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[10\].FF OVHB\[13\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[13\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07846__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11222_ _11216_/CLK line[49] VGND VGND VPWR VPWR _11222_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06172__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[7\].FF OVHB\[3\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[3\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[1\].TOBUF OVHB\[13\].VALID\[1\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12902__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11153_ _11152_/Q _11172_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10104_ _10100_/CLK line[50] VGND VGND VPWR VPWR _10105_/A sky130_fd_sc_hd__dfxtp_1
X_11084_ _11090_/CLK line[114] VGND VGND VPWR VPWR _11084_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11518__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10035_ _10034_/Q _10052_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08099__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[18\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11986_ _12002_/CLK line[29] VGND VGND VPWR VPWR _11986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13725_ _13725_/CLK _13726_/X VGND VGND VPWR VPWR _13701_/CLK sky130_fd_sc_hd__dlclkp_1
X_10937_ _10936_/Q _10962_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11253__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06347__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ _13907_/X wr VGND VGND VPWR VPWR _13656_/X sky130_fd_sc_hd__and2_1
XMUX.MUX\[9\] _11414_/Z _12884_/Z _13514_/Z _06864_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[9] sky130_fd_sc_hd__mux4_1
XANTENNA__05251__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10868_ _10872_/CLK line[30] VGND VGND VPWR VPWR _10868_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12607_ _12712_/A VGND VGND VPWR VPWR _12607_/Y sky130_fd_sc_hd__inv_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _13552_/A VGND VGND VPWR VPWR _13587_/Y sky130_fd_sc_hd__inv_2
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10799_ _10799_/A _10822_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08562__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12538_ _12560_/CLK line[16] VGND VGND VPWR VPWR _12538_/Q sky130_fd_sc_hd__dfxtp_1
X_12469_ _12468_/Q _12502_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].V OVHB\[29\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[29\].V/Q sky130_fd_sc_hd__dfrtp_1
XOVHB\[31\].VALID\[1\].FF OVHB\[31\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[31\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07178__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05010_ _05010_/CLK _05011_/X VGND VGND VPWR VPWR _05000_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06810__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06961_ _06960_/Q _06972_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11428__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08700_ _08710_/CLK line[63] VGND VGND VPWR VPWR _08700_/Q sky130_fd_sc_hd__dfxtp_1
X_05912_ _05902_/CLK line[54] VGND VGND VPWR VPWR _05912_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VOBUF OVHB\[16\].V/Q OVHB\[16\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_09680_ _09694_/CLK line[127] VGND VGND VPWR VPWR _09680_/Q sky130_fd_sc_hd__dfxtp_1
X_06892_ _06892_/CLK line[118] VGND VGND VPWR VPWR _06892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05426__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[1\].VALID\[9\].FF OVHB\[1\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[1\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08631_ _08630_/Q _08652_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_05843_ _05843_/A _05852_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13643__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[30\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08562_ _08560_/CLK line[113] VGND VGND VPWR VPWR _08562_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08737__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05774_ _05756_/CLK line[119] VGND VGND VPWR VPWR _05774_/Q sky130_fd_sc_hd__dfxtp_1
X_07513_ _07512_/Q _07532_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08493_ _08492_/Q _08512_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07444_ _07446_/CLK line[114] VGND VGND VPWR VPWR _07444_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05161__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09211__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07375_ _07374_/Q _07392_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09114_ _09116_/CLK line[124] VGND VGND VPWR VPWR _09114_/Q sky130_fd_sc_hd__dfxtp_1
X_06326_ _06320_/CLK line[115] VGND VGND VPWR VPWR _06327_/A sky130_fd_sc_hd__dfxtp_1
X_09045_ _09044_/Q _09072_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_06257_ _06256_/Q _06272_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12572__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07088__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05208_ _05214_/CLK line[116] VGND VGND VPWR VPWR _05209_/A sky130_fd_sc_hd__dfxtp_1
X_06188_ _06186_/CLK line[52] VGND VGND VPWR VPWR _06188_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12291__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13818__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05139_ _05139_/A _05152_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[12\].FF OVHB\[8\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[8\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05186__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09947_ _09912_/A VGND VGND VPWR VPWR _09947_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10242__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09878_ _09908_/CLK line[80] VGND VGND VPWR VPWR _09878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05336__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08829_ _08829_/A _08862_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13553__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11840_ _11846_/CLK line[90] VGND VGND VPWR VPWR _11840_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07551__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12169__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11771_ _11770_/Q _11802_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12747__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[6\].TOBUF OVHB\[11\].VALID\[6\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_13510_ _13509_/Q _13517_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10722_ _10728_/CLK line[91] VGND VGND VPWR VPWR _10722_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12466__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13441_ _13439_/CLK line[40] VGND VGND VPWR VPWR _13441_/Q sky130_fd_sc_hd__dfxtp_1
X_10653_ _10652_/Q _10682_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09478__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13372_ _13371_/Q _13377_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_10584_ _10594_/CLK line[28] VGND VGND VPWR VPWR _10584_/Q sky130_fd_sc_hd__dfxtp_1
X_12323_ _12311_/CLK line[41] VGND VGND VPWR VPWR _12324_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10417__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12254_ _12253_/Q _12257_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13728__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11205_ _11205_/CLK _11206_/X VGND VGND VPWR VPWR _11191_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12632__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _12185_/CLK _12186_/X VGND VGND VPWR VPWR _12177_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07726__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[4\].FF OVHB\[28\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[28\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11136_ _11311_/A wr VGND VGND VPWR VPWR _11136_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[4\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11067_ _11032_/A VGND VGND VPWR VPWR _11067_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09941__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10018_ _10042_/CLK line[16] VGND VGND VPWR VPWR _10018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[10\].VALID\[1\].FF OVHB\[10\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[10\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11969_ _11945_/CLK line[7] VGND VGND VPWR VPWR _11970_/A sky130_fd_sc_hd__dfxtp_1
X_13708_ _13708_/A _13727_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06077__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05490_ _05476_/CLK line[117] VGND VGND VPWR VPWR _05490_/Q sky130_fd_sc_hd__dfxtp_1
X_13639_ _13631_/CLK line[2] VGND VGND VPWR VPWR _13639_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12807__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[16\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09388__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08292__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07160_ _07170_/CLK line[127] VGND VGND VPWR VPWR _07160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06111_ _06110_/Q _06132_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_07091_ _07091_/A _07112_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06042_ _06050_/CLK line[113] VGND VGND VPWR VPWR _06042_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[12\].TOBUF OVHB\[16\].VALID\[12\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12542__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09801_ _09793_/CLK line[40] VGND VGND VPWR VPWR _09801_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06540__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07993_ _07992_/Q _08022_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11158__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09732_ _09731_/Q _09737_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_06944_ _06960_/CLK line[28] VGND VGND VPWR VPWR _06944_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09851__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[9\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09663_ _09659_/CLK line[105] VGND VGND VPWR VPWR _09664_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06875_ _06874_/Q _06902_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13373__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08614_ _08614_/A _08617_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08467__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05826_ _05836_/CLK line[29] VGND VGND VPWR VPWR _05827_/A sky130_fd_sc_hd__dfxtp_1
X_09594_ _09593_/Q _09597_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[26\].VALID\[6\].FF OVHB\[26\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[26\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08545_/CLK _08546_/X VGND VGND VPWR VPWR _08541_/CLK sky130_fd_sc_hd__dlclkp_1
X_05757_ _05757_/A _05782_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08476_ _13921_/X wr VGND VGND VPWR VPWR _08476_/X sky130_fd_sc_hd__and2_1
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05688_ _05708_/CLK line[94] VGND VGND VPWR VPWR _05688_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12717__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07427_ _13918_/X VGND VGND VPWR VPWR _07427_/Y sky130_fd_sc_hd__inv_2
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10087__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11621__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06715__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09876__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07358_ _07380_/CLK line[80] VGND VGND VPWR VPWR _07358_/Q sky130_fd_sc_hd__dfxtp_1
X_06309_ _06308_/Q _06342_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
X_07289_ _07288_/Q _07322_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_09028_ _09028_/A _09037_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13548__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[14\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06450__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11068__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13990_ _13990_/A _13990_/B _13982_/X _13990_/D VGND VGND VPWR VPWR _13990_/X sky130_fd_sc_hd__and4_4
XANTENNA__05066__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ _12937_/CLK line[67] VGND VGND VPWR VPWR _12941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13283__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08377__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _12871_/Q _12887_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07281__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[7\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _13270_/CLK sky130_fd_sc_hd__clkbuf_4
X_11823_ _11823_/CLK line[68] VGND VGND VPWR VPWR _11823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11381__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[0\].TOBUF OVHB\[26\].VALID\[0\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_11754_ _11754_/A _11767_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10707_/CLK line[69] VGND VGND VPWR VPWR _10705_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11691_/CLK line[5] VGND VGND VPWR VPWR _11685_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11531__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[8\].FF OVHB\[24\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[24\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13424_ _13423_/Q _13447_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_10636_ _10636_/A _10647_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06625__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[10\].FF OVHB\[4\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[4\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10147__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13355_ _13347_/CLK line[15] VGND VGND VPWR VPWR _13355_/Q sky130_fd_sc_hd__dfxtp_1
X_10567_ _10571_/CLK line[6] VGND VGND VPWR VPWR _10568_/A sky130_fd_sc_hd__dfxtp_1
X_12306_ _12306_/A _12327_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08840__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13286_ _13286_/A _13307_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_10498_ _10498_/A _10507_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13458__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12237_ _12227_/CLK line[1] VGND VGND VPWR VPWR _12237_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07456__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12168_ _12168_/A _12187_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11556__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11119_ _11111_/CLK line[2] VGND VGND VPWR VPWR _11119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12099_ _12109_/CLK line[66] VGND VGND VPWR VPWR _12100_/A sky130_fd_sc_hd__dfxtp_1
X_04990_ _05000_/CLK line[31] VGND VGND VPWR VPWR _04990_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].CGAND _09632_/A wr VGND VGND VPWR VPWR OVHB\[24\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11706__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06660_ _06682_/CLK line[26] VGND VGND VPWR VPWR _06660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07191__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05704__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05611_ _05610_/Q _05642_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_06591_ _06590_/Q _06622_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_08330_ _08329_/Q _08337_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_05542_ _05568_/CLK line[27] VGND VGND VPWR VPWR _05542_/Q sky130_fd_sc_hd__dfxtp_1
X_08261_ _08257_/CLK line[104] VGND VGND VPWR VPWR _08261_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[6\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _12885_/CLK sky130_fd_sc_hd__clkbuf_4
X_05473_ _05472_/Q _05502_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04928__A2_N _04918_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07212_ _07211_/Q _07217_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[6\].TOBUF OVHB\[18\].VALID\[6\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_08192_ _08192_/A _08197_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10057__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07143_ _07117_/CLK line[105] VGND VGND VPWR VPWR _07143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07074_ _07074_/A _07077_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[14\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06025_ _06025_/CLK _06026_/X VGND VGND VPWR VPWR _06023_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12272__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07366__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[1\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07976_ _07975_/Q _07987_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09581__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09715_ _09721_/CLK line[15] VGND VGND VPWR VPWR _09715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06927_ _06923_/CLK line[6] VGND VGND VPWR VPWR _06927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10520__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09646_ _09646_/A _09667_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _10225_/CLK sky130_fd_sc_hd__clkbuf_4
X_06858_ _06857_/Q _06867_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05614__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05809_ _05799_/CLK line[7] VGND VGND VPWR VPWR _05810_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09577_ _09577_/CLK line[65] VGND VGND VPWR VPWR _09578_/A sky130_fd_sc_hd__dfxtp_1
X_06789_ _06775_/CLK line[71] VGND VGND VPWR VPWR _06789_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08527_/Q _08547_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[18\].VALID\[10\].FF OVHB\[18\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[18\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12447__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _08473_/CLK line[66] VGND VGND VPWR VPWR _08459_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[27\] _10863_/Z _10373_/Z _11003_/Z _13593_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[27] sky130_fd_sc_hd__mux4_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ _11469_/Q _11487_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10421_ _10405_/CLK line[67] VGND VGND VPWR VPWR _10421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09756__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _13139_/Q _13167_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_10352_ _10352_/A _10367_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[0\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13071_ _13075_/CLK line[13] VGND VGND VPWR VPWR _13071_/Q sky130_fd_sc_hd__dfxtp_1
X_10283_ _10277_/CLK line[4] VGND VGND VPWR VPWR _10283_/Q sky130_fd_sc_hd__dfxtp_1
X_12022_ _12022_/A _12047_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06180__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[24\].VALID\[5\].TOBUF OVHB\[24\].VALID\[5\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12910__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13973_ _13979_/C _13979_/B _13979_/A _13979_/D VGND VGND VPWR VPWR _13973_/X sky130_fd_sc_hd__and4bb_4
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12924_ _12923_/Q _12957_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12855_ _12881_/CLK line[42] VGND VGND VPWR VPWR _12855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11806_ _11805_/Q _11837_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_12786_ _12785_/Q _12817_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[25\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _09840_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _11757_/CLK line[43] VGND VGND VPWR VPWR _11737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11261__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].CGAND_A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06355__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _11667_/Q _11697_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13406_/Q _13412_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_10619_ _10627_/CLK line[44] VGND VGND VPWR VPWR _10619_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11599_ _11605_/CLK line[108] VGND VGND VPWR VPWR _11600_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08570__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13338_ _13308_/CLK line[121] VGND VGND VPWR VPWR _13339_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13188__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13269_ _13268_/Q _13272_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07830_ _07829_/Q _07847_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12820__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07761_ _07773_/CLK line[3] VGND VGND VPWR VPWR _07761_/Q sky130_fd_sc_hd__dfxtp_1
X_04973_ _04947_/CLK line[9] VGND VGND VPWR VPWR _04973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11436__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09500_ _09499_/Q _09527_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[15\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06712_ _06712_/A _06727_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_07692_ _07691_/Q _07707_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09431_ _09427_/CLK line[13] VGND VGND VPWR VPWR _09431_/Q sky130_fd_sc_hd__dfxtp_1
X_06643_ _06633_/CLK line[4] VGND VGND VPWR VPWR _06643_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[4\].TOBUF OVHB\[30\].VALID\[4\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13651__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09362_ _09361_/Q _09387_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08745__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06574_ _06573_/Q _06587_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_08313_ _08329_/CLK line[14] VGND VGND VPWR VPWR _08313_/Q sky130_fd_sc_hd__dfxtp_1
X_05525_ _05519_/CLK line[5] VGND VGND VPWR VPWR _05525_/Q sky130_fd_sc_hd__dfxtp_1
X_09293_ _09307_/CLK line[78] VGND VGND VPWR VPWR _09293_/Q sky130_fd_sc_hd__dfxtp_1
X_08244_ _08244_/A _08267_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05456_ _05455_/Q _05467_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08175_ _08175_/CLK line[79] VGND VGND VPWR VPWR _08176_/A sky130_fd_sc_hd__dfxtp_1
X_05387_ _05391_/CLK line[70] VGND VGND VPWR VPWR _05387_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _09455_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[28\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07126_ _07125_/Q _07147_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08480__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13098__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[14\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _06585_/CLK sky130_fd_sc_hd__clkbuf_4
X_07057_ _07043_/CLK line[65] VGND VGND VPWR VPWR _07057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07096__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06008_ _06007_/Q _06027_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13826__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07959_ _07981_/CLK line[108] VGND VGND VPWR VPWR _07960_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DEC.DEC0.AND1_A_N A[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10250__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].CG clk OVHB\[14\].CGAND/X VGND VGND VPWR VPWR OVHB\[14\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10970_ _10970_/A _10997_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05344__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05922__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09629_ _09629_/A _09632_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13561__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05641__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _12640_/CLK _12641_/X VGND VGND VPWR VPWR _12638_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08655__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12177__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _12712_/A wr VGND VGND VPWR VPWR _12571_/X sky130_fd_sc_hd__and2_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _11592_/A VGND VGND VPWR VPWR _11522_/Y sky130_fd_sc_hd__inv_2
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _11479_/CLK line[32] VGND VGND VPWR VPWR _11453_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[6\].VALID\[14\].TOBUF OVHB\[6\].VALID\[14\].FF/Q OVHB\[6\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__09486__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10404_ _10403_/Q _10437_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06903__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11384_ _11383_/Q _11417_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13586__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13123_ _13123_/A _13132_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_10335_ _10341_/CLK line[42] VGND VGND VPWR VPWR _10335_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10425__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[1\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05519__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _13050_/CLK line[119] VGND VGND VPWR VPWR _13054_/Q sky130_fd_sc_hd__dfxtp_1
X_10266_ _10265_/Q _10297_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13736__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12005_ _12004_/Q _12012_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05816__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10197_ _10217_/CLK line[107] VGND VGND VPWR VPWR _10197_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[13\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _06200_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_79_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07734__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10160__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[27\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13956_ _13950_/A _13950_/B _13950_/C _13957_/D VGND VGND VPWR VPWR _13956_/X sky130_fd_sc_hd__and4b_4
XFILLER_46_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[19\]_A3 _07167_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12907_ _12906_/Q _12922_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_13887_ _13886_/Q _13902_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12838_ _12820_/CLK line[20] VGND VGND VPWR VPWR _12839_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[10\].TOBUF OVHB\[26\].VALID\[10\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_50_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12087__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _12769_/A _12782_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_05310_ _05309_/Q _05327_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06085__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06290_ _06290_/A _06307_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05241_ _05253_/CLK line[3] VGND VGND VPWR VPWR _05242_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07909__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09396__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05172_ _05171_/Q _05187_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[19\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10335__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09980_ _09980_/CLK _09981_/X VGND VGND VPWR VPWR _09978_/CLK sky130_fd_sc_hd__dlclkp_1
X_08931_ _13923_/X wr VGND VGND VPWR VPWR _08931_/X sky130_fd_sc_hd__and2_1
XOVHB\[6\].VALID\[2\].TOBUF OVHB\[6\].VALID\[2\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12550__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08862_ _13922_/X VGND VGND VPWR VPWR _08862_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07644__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07813_ _07837_/CLK line[32] VGND VGND VPWR VPWR _07813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08793_ _08823_/CLK line[96] VGND VGND VPWR VPWR _08793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11166__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07744_ _07743_/Q _07777_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04956_ _04955_/Q _04977_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[12\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _05815_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07675_ _07679_/CLK line[106] VGND VGND VPWR VPWR _07675_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].CG clk OVHB\[9\].CGAND/X VGND VGND VPWR VPWR OVHB\[9\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09414_ _09414_/CLK line[119] VGND VGND VPWR VPWR _09414_/Q sky130_fd_sc_hd__dfxtp_1
X_06626_ _06625_/Q _06657_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_MUX.MUX\[1\]_A1 _13428_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09345_ _09344_/Q _09352_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_06557_ _06565_/CLK line[107] VGND VGND VPWR VPWR _06558_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05508_ _05508_/A _05537_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
X_09276_ _09256_/CLK line[56] VGND VGND VPWR VPWR _09277_/A sky130_fd_sc_hd__dfxtp_1
X_06488_ _06487_/Q _06517_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_08227_ _08226_/Q _08232_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12725__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05439_ _05445_/CLK line[108] VGND VGND VPWR VPWR _05439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07819__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06723__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08158_ _08134_/CLK line[57] VGND VGND VPWR VPWR _08158_/Q sky130_fd_sc_hd__dfxtp_1
X_07109_ _07109_/A _07112_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_08089_ _08088_/Q _08092_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10120_ _10120_/CLK _10121_/X VGND VGND VPWR VPWR _10100_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[26\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10051_ _10192_/A wr VGND VGND VPWR VPWR _10051_/X sky130_fd_sc_hd__and2_1
XFILLER_130_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11076__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _13822_/CLK line[95] VGND VGND VPWR VPWR _13810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05074__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13741_ _13741_/A _13762_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_10953_ _10952_/Q _10962_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13291__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[10\].FF OVHB\[9\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[9\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08385__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13672_ _13682_/CLK line[17] VGND VGND VPWR VPWR _13672_/Q sky130_fd_sc_hd__dfxtp_1
X_10884_ _10872_/CLK line[23] VGND VGND VPWR VPWR _10885_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ _12623_/A _12642_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _12560_/CLK line[18] VGND VGND VPWR VPWR _12554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11505_/A _11522_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ _12484_/Q _12502_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06633__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11436_ _11440_/CLK line[19] VGND VGND VPWR VPWR _11436_/Q sky130_fd_sc_hd__dfxtp_1
X_11367_ _11367_/A _11382_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05249__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13106_ _13120_/CLK line[29] VGND VGND VPWR VPWR _13106_/Q sky130_fd_sc_hd__dfxtp_1
X_10318_ _10314_/CLK line[20] VGND VGND VPWR VPWR _10319_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11298_ _11302_/CLK line[84] VGND VGND VPWR VPWR _11298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13466__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13037_ _13036_/Q _13062_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_10249_ _10249_/A _10262_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05790_ _05789_/Q _05817_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13939_ _13944_/B _13946_/B _13944_/C _13944_/D VGND VGND VPWR VPWR _05152_/A sky130_fd_sc_hd__nor4b_4
XANTENNA__11714__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06808__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07460_ _07460_/CLK _07461_/X VGND VGND VPWR VPWR _07446_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_50_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06411_ _06551_/A wr VGND VGND VPWR VPWR _06411_/X sky130_fd_sc_hd__and2_1
X_07391_ _13918_/X wr VGND VGND VPWR VPWR _07391_/X sky130_fd_sc_hd__and2_1
XFILLER_124_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09130_ _09116_/CLK line[117] VGND VGND VPWR VPWR _09131_/A sky130_fd_sc_hd__dfxtp_1
X_06342_ _06272_/A VGND VGND VPWR VPWR _06342_/Y sky130_fd_sc_hd__inv_2
XOVHB\[4\].VALID\[7\].TOBUF OVHB\[4\].VALID\[7\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VOBUF OVHB\[12\].V/Q OVHB\[12\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_09061_ _09061_/A _09072_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_06273_ _06285_/CLK line[96] VGND VGND VPWR VPWR _06273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08012_ _08000_/CLK line[118] VGND VGND VPWR VPWR _08012_/Q sky130_fd_sc_hd__dfxtp_1
X_05224_ _05224_/A _05257_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10065__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05155_ _05157_/CLK line[106] VGND VGND VPWR VPWR _05155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05159__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09963_ _09962_/Q _09982_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_05086_ _05085_/Q _05117_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12280__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08914_ _08922_/CLK line[18] VGND VGND VPWR VPWR _08914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__04998__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09894_ _09908_/CLK line[82] VGND VGND VPWR VPWR _09894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07374__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07952__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08845_ _08845_/A _08862_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07671__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08776_ _08762_/CLK line[83] VGND VGND VPWR VPWR _08776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05988_ _05984_/CLK line[89] VGND VGND VPWR VPWR _05988_/Q sky130_fd_sc_hd__dfxtp_1
X_07727_ _07726_/Q _07742_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_04939_ A_h[13] _04939_/B2 A_h[13] _04939_/B2 VGND VGND VPWR VPWR _04941_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07658_ _07644_/CLK line[84] VGND VGND VPWR VPWR _07658_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05622__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[20\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06609_ _06608_/Q _06622_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_07589_ _07589_/A _07602_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09328_ _09320_/CLK line[94] VGND VGND VPWR VPWR _09328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08933__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[9\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[19\].VALID\[0\].FF OVHB\[19\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[19\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12455__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09259_ _09258_/Q _09282_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07549__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12270_ _12268_/CLK line[31] VGND VGND VPWR VPWR _12270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11221_ _11220_/Q _11242_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07846__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09764__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11152_ _11148_/CLK line[17] VGND VGND VPWR VPWR _11152_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[2\].TOBUF OVHB\[11\].VALID\[2\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_62_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10103_ _10102_/Q _10122_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12190__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10703__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11083_ _11082_/Q _11102_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_10034_ _10042_/CLK line[18] VGND VGND VPWR VPWR _10034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[17\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[24\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _11985_/A _12012_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13724_ _13724_/A _13727_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_10936_ _10930_/CLK line[61] VGND VGND VPWR VPWR _10936_/Q sky130_fd_sc_hd__dfxtp_1
X_13655_ _13655_/CLK _13656_/X VGND VGND VPWR VPWR _13631_/CLK sky130_fd_sc_hd__dlclkp_1
X_10867_ _10866_/Q _10892_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09939__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12712_/A wr VGND VGND VPWR VPWR _12606_/X sky130_fd_sc_hd__and2_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ _13552_/A wr VGND VGND VPWR VPWR _13586_/X sky130_fd_sc_hd__and2_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ _10804_/CLK line[126] VGND VGND VPWR VPWR _10799_/A sky130_fd_sc_hd__dfxtp_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12365__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12537_ _12712_/A VGND VGND VPWR VPWR _12537_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06363__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12468_ _12490_/CLK line[112] VGND VGND VPWR VPWR _12468_/Q sky130_fd_sc_hd__dfxtp_1
X_11419_ _11419_/A _11452_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_12399_ _12398_/Q _12432_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09674__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[2\].FF OVHB\[17\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[17\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13196__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[4\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _12500_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10613__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06960_ _06960_/CLK line[21] VGND VGND VPWR VPWR _06960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05911_ _05911_/A _05922_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_06891_ _06891_/A _06902_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_08630_ _08646_/CLK line[31] VGND VGND VPWR VPWR _08630_/Q sky130_fd_sc_hd__dfxtp_1
X_05842_ _05836_/CLK line[22] VGND VGND VPWR VPWR _05843_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07922__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05292__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08561_ _08560_/Q _08582_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_05773_ _05772_/Q _05782_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11444__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07512_ _07518_/CLK line[17] VGND VGND VPWR VPWR _07512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06538__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08492_ _08480_/CLK line[81] VGND VGND VPWR VPWR _08492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07443_ _07443_/A _07462_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09849__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08753__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07374_ _07380_/CLK line[82] VGND VGND VPWR VPWR _07374_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09211__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09113_ _09113_/A _09142_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
X_06325_ _06324_/Q _06342_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13949__A A_h[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].CGAND _13920_/X wr VGND VGND VPWR VPWR OVHB\[19\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__06273__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09044_ _09068_/CLK line[92] VGND VGND VPWR VPWR _09044_/Q sky130_fd_sc_hd__dfxtp_1
X_06256_ _06244_/CLK line[83] VGND VGND VPWR VPWR _06256_/Q sky130_fd_sc_hd__dfxtp_1
X_05207_ _05206_/Q _05222_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06187_ _06186_/Q _06202_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05467__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05138_ _05122_/CLK line[84] VGND VGND VPWR VPWR _05139_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11619__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05186__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09946_ _09912_/A wr VGND VGND VPWR VPWR _09946_/X sky130_fd_sc_hd__and2_1
X_05069_ _05068_/Q _05082_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09877_ _09912_/A VGND VGND VPWR VPWR _09877_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[3\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _12115_/CLK sky130_fd_sc_hd__clkbuf_4
X_08828_ _08850_/CLK line[112] VGND VGND VPWR VPWR _08829_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08928__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[4\].FF OVHB\[15\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[15\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ _08759_/A _08792_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11354__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06448__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ _11776_/CLK line[58] VGND VGND VPWR VPWR _11770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05352__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10721_ _10720_/Q _10752_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[13\].FF OVHB\[31\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[31\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13440_ _13439_/Q _13447_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08663__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10652_ _10656_/CLK line[59] VGND VGND VPWR VPWR _10652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13371_ _13347_/CLK line[8] VGND VGND VPWR VPWR _13371_/Q sky130_fd_sc_hd__dfxtp_1
X_10583_ _10583_/A _10612_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07279__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _12321_/Q _12327_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06761__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12253_ _12227_/CLK line[9] VGND VGND VPWR VPWR _12253_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[14\].TOBUF OVHB\[19\].VALID\[14\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_11204_ _11204_/A _11207_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06911__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12184_ _12184_/A _12187_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11529__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11135_ _11135_/CLK _11136_/X VGND VGND VPWR VPWR _11111_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10433__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05527__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11066_ _11032_/A wr VGND VGND VPWR VPWR _11066_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[17\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13744__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10017_ _10192_/A VGND VGND VPWR VPWR _10017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08838__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11968_ _11967_/Q _11977_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06936__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05262__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[2\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _11170_/CLK sky130_fd_sc_hd__clkbuf_4
X_13707_ _13701_/CLK line[33] VGND VGND VPWR VPWR _13708_/A sky130_fd_sc_hd__dfxtp_1
X_10919_ _10903_/CLK line[39] VGND VGND VPWR VPWR _10919_/Q sky130_fd_sc_hd__dfxtp_1
X_11899_ _11901_/CLK line[103] VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[13\].VALID\[6\].FF OVHB\[13\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[13\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[13\].TOBUF OVHB\[12\].VALID\[13\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_13638_ _13638_/A _13657_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[27\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[22\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12095__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10608__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].CGAND _13921_/X wr VGND VGND VPWR VPWR OVHB\[20\].CG/GATE sky130_fd_sc_hd__and2_4
XFILLER_30_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13569_ _13559_/CLK line[98] VGND VGND VPWR VPWR _13569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07189__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06110_ _06108_/CLK line[31] VGND VGND VPWR VPWR _06110_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06093__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07090_ _07098_/CLK line[95] VGND VGND VPWR VPWR _07091_/A sky130_fd_sc_hd__dfxtp_1
X_06041_ _06040_/Q _06062_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09982__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10343__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09800_ _09799_/Q _09807_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07992_ _08000_/CLK line[123] VGND VGND VPWR VPWR _07992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05437__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09731_ _09721_/CLK line[8] VGND VGND VPWR VPWR _09731_/Q sky130_fd_sc_hd__dfxtp_1
X_06943_ _06942_/Q _06972_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[2\].TOBUF OVHB\[18\].VALID\[2\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_80_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[22\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _09070_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09662_ _09661_/Q _09667_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06874_ _06892_/CLK line[124] VGND VGND VPWR VPWR _06874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07652__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08613_ _08609_/CLK line[9] VGND VGND VPWR VPWR _08614_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07007__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05825_ _05824_/Q _05852_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_09593_ _09577_/CLK line[73] VGND VGND VPWR VPWR _09593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _08544_/A _08547_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06268__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05756_ _05756_/CLK line[125] VGND VGND VPWR VPWR _05757_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _08475_/CLK _08476_/X VGND VGND VPWR VPWR _08473_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05687_ _05687_/A _05712_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09579__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07426_ _13918_/X wr VGND VGND VPWR VPWR _07426_/X sky130_fd_sc_hd__and2_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05900__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07357_ _13918_/X VGND VGND VPWR VPWR _07357_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10518__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09876__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06308_ _06320_/CLK line[112] VGND VGND VPWR VPWR _06308_/Q sky130_fd_sc_hd__dfxtp_1
X_07288_ _07292_/CLK line[48] VGND VGND VPWR VPWR _07288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09027_ _09005_/CLK line[70] VGND VGND VPWR VPWR _09028_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12733__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06239_ _06238_/Q _06272_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[20\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[8\].FF OVHB\[11\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[11\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07827__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09929_ _09925_/CLK line[98] VGND VGND VPWR VPWR _09929_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08301__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12940_ _12939_/Q _12957_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12871_ _12881_/CLK line[35] VGND VGND VPWR VPWR _12871_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11084__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11662__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06178__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ _11821_/Q _11837_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[21\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _08685_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11381__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11753_ _11757_/CLK line[36] VGND VGND VPWR VPWR _11754_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12908__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[24\].VALID\[1\].TOBUF OVHB\[24\].VALID\[1\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10703_/Q _10717_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08393__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11684_/A _11697_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _10627_/CLK line[37] VGND VGND VPWR VPWR _10636_/A sky130_fd_sc_hd__dfxtp_1
X_13423_ _13439_/CLK line[46] VGND VGND VPWR VPWR _13423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13354_ _13353_/Q _13377_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_10566_ _10565_/Q _10577_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_12305_ _12311_/CLK line[47] VGND VGND VPWR VPWR _12306_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12643__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13285_ _13285_/CLK line[111] VGND VGND VPWR VPWR _13286_/A sky130_fd_sc_hd__dfxtp_1
X_10497_ _10473_/CLK line[102] VGND VGND VPWR VPWR _10498_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12236_ _12236_/A _12257_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06641__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11259__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11837__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12167_ _12177_/CLK line[97] VGND VGND VPWR VPWR _12168_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09952__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11118_ _11118_/A _11137_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11556__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12098_/A _12117_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13474__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11049_ _11063_/CLK line[98] VGND VGND VPWR VPWR _11050_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08568__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05610_ _05632_/CLK line[58] VGND VGND VPWR VPWR _05610_/Q sky130_fd_sc_hd__dfxtp_1
X_06590_ _06596_/CLK line[122] VGND VGND VPWR VPWR _06590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05541_ _05541_/A _05572_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12818__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11722__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08260_ _08259_/Q _08267_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06816__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05472_ _05476_/CLK line[123] VGND VGND VPWR VPWR _05472_/Q sky130_fd_sc_hd__dfxtp_1
X_07211_ _07183_/CLK line[8] VGND VGND VPWR VPWR _07211_/Q sky130_fd_sc_hd__dfxtp_1
X_08191_ _08175_/CLK line[72] VGND VGND VPWR VPWR _08192_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[7\].TOBUF OVHB\[16\].VALID\[7\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_07142_ _07141_/Q _07147_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07497__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _05430_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13649__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07073_ _07043_/CLK line[73] VGND VGND VPWR VPWR _07074_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06024_ _06023_/Q _06027_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[0\].TOBUF OVHB\[30\].VALID\[0\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10073__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05167__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07975_ _07981_/CLK line[101] VGND VGND VPWR VPWR _07975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13384__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09714_ _09714_/A _09737_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_06926_ _06925_/Q _06937_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08478__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07382__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09645_ _09659_/CLK line[111] VGND VGND VPWR VPWR _09646_/A sky130_fd_sc_hd__dfxtp_1
X_06857_ _06839_/CLK line[102] VGND VGND VPWR VPWR _06857_/Q sky130_fd_sc_hd__dfxtp_1
X_05808_ _05807_/Q _05817_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09576_ _09575_/Q _09597_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06788_ _06788_/A _06797_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08541_/CLK line[97] VGND VGND VPWR VPWR _08527_/Q sky130_fd_sc_hd__dfxtp_1
X_05739_ _05739_/CLK line[103] VGND VGND VPWR VPWR _05740_/A sky130_fd_sc_hd__dfxtp_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _08457_/Q _08477_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05630__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07393_/CLK line[98] VGND VGND VPWR VPWR _07410_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10248__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08389_ _08383_/CLK line[34] VGND VGND VPWR VPWR _08389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13202__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10420_ _10419_/Q _10437_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08941__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13559__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10351_ _10341_/CLK line[35] VGND VGND VPWR VPWR _10352_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12463__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07557__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13070_ _13069_/Q _13097_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_10282_ _10281_/Q _10297_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[4\].VALID\[1\].FF OVHB\[4\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[4\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12021_ _12019_/CLK line[45] VGND VGND VPWR VPWR _12022_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[6\].TOBUF OVHB\[22\].VALID\[6\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11807__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10711__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13972_ _13979_/A _13979_/B _13979_/C _13979_/D VGND VGND VPWR VPWR _13972_/Y sky130_fd_sc_hd__nor4b_4
XANTENNA__08966__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07292__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05805__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12923_ _12937_/CLK line[64] VGND VGND VPWR VPWR _12923_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[10\].TOBUF OVHB\[6\].VALID\[10\].FF/Q OVHB\[6\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_100_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12854_ _12853_/Q _12887_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[7\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12638__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11805_ _11823_/CLK line[74] VGND VGND VPWR VPWR _11805_/Q sky130_fd_sc_hd__dfxtp_1
X_12785_ _12803_/CLK line[10] VGND VGND VPWR VPWR _12785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11736_ _11735_/Q _11767_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05540__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10158__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ _11691_/CLK line[11] VGND VGND VPWR VPWR _11667_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13394_/CLK line[24] VGND VGND VPWR VPWR _13406_/Q sky130_fd_sc_hd__dfxtp_1
X_10618_ _10617_/Q _10647_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _11597_/Q _11627_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[18\].CGAND_A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[18\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12373__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10549_ _10571_/CLK line[12] VGND VGND VPWR VPWR _10549_/Q sky130_fd_sc_hd__dfxtp_1
X_13337_ _13336_/Q _13342_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07467__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06371__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13254_/CLK line[89] VGND VGND VPWR VPWR _13268_/Q sky130_fd_sc_hd__dfxtp_1
X_12219_ _12218_/Q _12222_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[15\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _13198_/Q _13202_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10471__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09682__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09037__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10621__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07760_ _07759_/Q _07777_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08298__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04972_ _04971_/Q _04977_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05715__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06711_ _06711_/CLK line[35] VGND VGND VPWR VPWR _06712_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[3\].FF OVHB\[2\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[2\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07691_ _07679_/CLK line[99] VGND VGND VPWR VPWR _07691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09430_ _09429_/Q _09457_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_06642_ _06641_/Q _06657_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07930__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09361_ _09365_/CLK line[109] VGND VGND VPWR VPWR _09361_/Q sky130_fd_sc_hd__dfxtp_1
X_06573_ _06565_/CLK line[100] VGND VGND VPWR VPWR _06573_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12548__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08312_ _08311_/Q _08337_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_05524_ _05524_/A _05537_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06546__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09292_ _09291_/Q _09317_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[8\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08243_ _08257_/CLK line[110] VGND VGND VPWR VPWR _08244_/A sky130_fd_sc_hd__dfxtp_1
X_05455_ _05445_/CLK line[101] VGND VGND VPWR VPWR _05455_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10646__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09857__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _08173_/Q _08197_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05386_ _05385_/Q _05397_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07125_ _07117_/CLK line[111] VGND VGND VPWR VPWR _07125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06281__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07056_ _07056_/A _07077_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_06007_ _06023_/CLK line[97] VGND VGND VPWR VPWR _06007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13692__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07958_ _07958_/A _07987_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_06909_ _06923_/CLK line[12] VGND VGND VPWR VPWR _06909_/Q sky130_fd_sc_hd__dfxtp_1
X_07889_ _07905_/CLK line[76] VGND VGND VPWR VPWR _07889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09628_ _09626_/CLK line[89] VGND VGND VPWR VPWR _09629_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[29\].VALID\[12\].TOBUF OVHB\[29\].VALID\[12\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _09558_/Q _09562_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11362__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06456__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12570_ _12570_/CLK _12571_/X VGND VGND VPWR VPWR _12560_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[0\].VALID\[5\].FF OVHB\[0\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[0\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11592_/A wr VGND VGND VPWR VPWR _11521_/X sky130_fd_sc_hd__and2_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08671__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11452_ _11592_/A VGND VGND VPWR VPWR _11452_/Y sky130_fd_sc_hd__inv_2
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13289__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10403_ _10405_/CLK line[64] VGND VGND VPWR VPWR _10403_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13867__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11383_ _11395_/CLK line[0] VGND VGND VPWR VPWR _11383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10334_ _10333_/Q _10367_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_13122_ _13120_/CLK line[22] VGND VGND VPWR VPWR _13123_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13586__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13053_ _13052_/Q _13062_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_10265_ _10277_/CLK line[10] VGND VGND VPWR VPWR _10265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12004_ _12002_/CLK line[23] VGND VGND VPWR VPWR _12004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10196_ _10195_/Q _10227_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11537__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[22\].VALID\[11\].TOBUF OVHB\[22\].VALID\[11\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09007__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[27\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13955_ _13950_/B _13950_/A _13950_/C _13957_/D VGND VGND VPWR VPWR _13955_/X sky130_fd_sc_hd__and4b_4
XANTENNA__13752__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12906_ _12902_/CLK line[51] VGND VGND VPWR VPWR _12906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08846__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12011__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13886_ _13882_/CLK line[115] VGND VGND VPWR VPWR _13886_/Q sky130_fd_sc_hd__dfxtp_1
X_12837_ _12836_/Q _12852_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05270__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12768_ _12774_/CLK line[116] VGND VGND VPWR VPWR _12769_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11719_ _11719_/A _11732_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12699_ _12698_/Q _12712_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_05240_ _05239_/Q _05257_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05171_ _05157_/CLK line[99] VGND VGND VPWR VPWR _05171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07197__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08930_ _08930_/CLK _08931_/X VGND VGND VPWR VPWR _08922_/CLK sky130_fd_sc_hd__dlclkp_1
X_08861_ _13922_/X wr VGND VGND VPWR VPWR _08861_/X sky130_fd_sc_hd__and2_1
XFILLER_111_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10351__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[3\].TOBUF OVHB\[4\].VALID\[3\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_07812_ _13920_/X VGND VGND VPWR VPWR _07812_/Y sky130_fd_sc_hd__inv_2
X_08792_ _13922_/X VGND VGND VPWR VPWR _08792_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05445__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[2\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[6\].TOBUF OVHB\[29\].VALID\[6\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_07743_ _07773_/CLK line[0] VGND VGND VPWR VPWR _07743_/Q sky130_fd_sc_hd__dfxtp_1
X_04955_ _04947_/CLK line[15] VGND VGND VPWR VPWR _04955_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[13\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13662__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07674_ _07673_/Q _07707_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07660__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[0\].FF OVHB\[27\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[27\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06625_ _06633_/CLK line[10] VGND VGND VPWR VPWR _06625_/Q sky130_fd_sc_hd__dfxtp_1
X_09413_ _09412_/Q _09422_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12278__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[12\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[1\]_A2 _13498_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06556_ _06556_/A _06587_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_09344_ _09320_/CLK line[87] VGND VGND VPWR VPWR _09344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05507_ _05519_/CLK line[11] VGND VGND VPWR VPWR _05508_/A sky130_fd_sc_hd__dfxtp_1
X_09275_ _09274_/Q _09282_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_06487_ _06489_/CLK line[75] VGND VGND VPWR VPWR _06487_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11910__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09587__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08226_ _08208_/CLK line[88] VGND VGND VPWR VPWR _08226_/Q sky130_fd_sc_hd__dfxtp_1
X_05438_ _05438_/A _05467_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_08157_ _08156_/Q _08162_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10526__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05369_ _05391_/CLK line[76] VGND VGND VPWR VPWR _05369_/Q sky130_fd_sc_hd__dfxtp_1
X_07108_ _07098_/CLK line[89] VGND VGND VPWR VPWR _07109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[6\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08088_ _08070_/CLK line[25] VGND VGND VPWR VPWR _08088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13837__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12741__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07039_ _07038_/Q _07042_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07835__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10050_ _10050_/CLK _10051_/X VGND VGND VPWR VPWR _10042_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_88_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[31\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _11940_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[3\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13740_ _13746_/CLK line[63] VGND VGND VPWR VPWR _13741_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10952_ _10930_/CLK line[54] VGND VGND VPWR VPWR _10952_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07570__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12188__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13671_ _13670_/Q _13692_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11092__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10883_ _10882_/Q _10892_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06186__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ _12638_/CLK line[49] VGND VGND VPWR VPWR _12623_/A sky130_fd_sc_hd__dfxtp_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _12552_/Q _12572_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09497__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _11500_/CLK line[50] VGND VGND VPWR VPWR _11505_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[25\].VALID\[2\].FF OVHB\[25\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[25\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12490_/CLK line[114] VGND VGND VPWR VPWR _12484_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ _11434_/Q _11452_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _05185_/CLK sky130_fd_sc_hd__clkbuf_4
X_11366_ _11370_/CLK line[115] VGND VGND VPWR VPWR _11367_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12651__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13105_ _13104_/Q _13132_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_10317_ _10316_/Q _10332_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_11297_ _11297_/A _11312_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07745__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10248_ _10248_/CLK line[116] VGND VGND VPWR VPWR _10249_/A sky130_fd_sc_hd__dfxtp_1
X_13036_ _13050_/CLK line[125] VGND VGND VPWR VPWR _13036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11267__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10179_ _10178_/Q _10192_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09960__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08576__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13938_ A[6] VGND VGND VPWR VPWR _13944_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_OVHB\[25\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13869_ _13868_/Q _13902_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12676__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[30\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _11555_/CLK sky130_fd_sc_hd__clkbuf_4
X_06410_ _06410_/CLK _06411_/X VGND VGND VPWR VPWR _06408_/CLK sky130_fd_sc_hd__dlclkp_1
X_07390_ _07390_/CLK _07391_/X VGND VGND VPWR VPWR _07380_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_22_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06341_ _06272_/A wr VGND VGND VPWR VPWR _06341_/X sky130_fd_sc_hd__and2_1
XANTENNA__12826__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[13\].FF OVHB\[22\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[22\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[8\].TOBUF OVHB\[2\].VALID\[8\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_09060_ _09068_/CLK line[85] VGND VGND VPWR VPWR _09061_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06824__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06272_ _06272_/A VGND VGND VPWR VPWR _06272_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09200__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08011_ _08010_/Q _08022_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_05223_ _05253_/CLK line[0] VGND VGND VPWR VPWR _05224_/A sky130_fd_sc_hd__dfxtp_1
X_05154_ _05153_/Q _05187_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04922__A A_h[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09962_ _09978_/CLK line[113] VGND VGND VPWR VPWR _09962_/Q sky130_fd_sc_hd__dfxtp_1
X_05085_ _05093_/CLK line[74] VGND VGND VPWR VPWR _05085_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[4\].FF OVHB\[23\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[23\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08913_ _08912_/Q _08932_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_09893_ _09892_/Q _09912_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11177__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10081__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08844_ _08850_/CLK line[114] VGND VGND VPWR VPWR _08845_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05175__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].CGAND _06832_/A wr VGND VGND VPWR VPWR OVHB\[15\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_100_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05987_ _05986_/Q _05992_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_08775_ _08775_/A _08792_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13392__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13970__A A_h[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04938_ A_h[10] _04938_/B2 A_h[10] _04938_/B2 VGND VGND VPWR VPWR _04938_/X sky130_fd_sc_hd__a2bb2o_4
X_07726_ _07724_/CLK line[115] VGND VGND VPWR VPWR _07726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08486__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07657_ _07656_/Q _07672_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06608_ _06596_/CLK line[116] VGND VGND VPWR VPWR _06608_/Q sky130_fd_sc_hd__dfxtp_1
X_07588_ _07572_/CLK line[52] VGND VGND VPWR VPWR _07589_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[11\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06539_ _06538_/Q _06552_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_09327_ _09327_/A _09352_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_MUX.MUX\[9\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11640__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06734__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09258_ _09256_/CLK line[62] VGND VGND VPWR VPWR _09258_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09110__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10256__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08209_ _08209_/A _08232_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_09189_ _09188_/Q _09212_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[17\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11220_ _11216_/CLK line[63] VGND VGND VPWR VPWR _11220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13567__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ _11150_/Q _11172_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10102_ _10100_/CLK line[49] VGND VGND VPWR VPWR _10102_/Q sky130_fd_sc_hd__dfxtp_1
X_11082_ _11090_/CLK line[113] VGND VGND VPWR VPWR _11082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10033_ _10032_/Q _10052_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[4\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05085__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11815__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[6\].FF OVHB\[21\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[21\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06909__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05813__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11984_ _12002_/CLK line[28] VGND VGND VPWR VPWR _11985_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[30\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[19\].VALID\[10\].TOBUF OVHB\[19\].VALID\[10\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_13723_ _13701_/CLK line[41] VGND VGND VPWR VPWR _13724_/A sky130_fd_sc_hd__dfxtp_1
X_10935_ _10934_/Q _10962_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _13653_/Q _13657_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_10866_ _10872_/CLK line[29] VGND VGND VPWR VPWR _10866_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _12605_/CLK _12606_/X VGND VGND VPWR VPWR _12601_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _13585_/CLK _13586_/X VGND VGND VPWR VPWR _13559_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[27\].CG clk OVHB\[27\].CGAND/X VGND VGND VPWR VPWR OVHB\[27\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_10797_ _10796_/Q _10822_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12536_ _12712_/A wr VGND VGND VPWR VPWR _12536_/X sky130_fd_sc_hd__and2_1
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10166__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12467_ _13943_/X VGND VGND VPWR VPWR _12467_/Y sky130_fd_sc_hd__inv_2
X_11418_ _11440_/CLK line[16] VGND VGND VPWR VPWR _11419_/A sky130_fd_sc_hd__dfxtp_1
X_12398_ _12414_/CLK line[80] VGND VGND VPWR VPWR _12398_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12381__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11349_ _11348_/Q _11382_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07475__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05910_ _05902_/CLK line[53] VGND VGND VPWR VPWR _05911_/A sky130_fd_sc_hd__dfxtp_1
X_13019_ _12999_/CLK line[103] VGND VGND VPWR VPWR _13019_/Q sky130_fd_sc_hd__dfxtp_1
X_06890_ _06892_/CLK line[117] VGND VGND VPWR VPWR _06891_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09690__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05841_ _05841_/A _05852_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_08560_ _08560_/CLK line[127] VGND VGND VPWR VPWR _08560_/Q sky130_fd_sc_hd__dfxtp_1
X_05772_ _05756_/CLK line[118] VGND VGND VPWR VPWR _05772_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05723__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07511_ _07510_/Q _07532_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
X_08491_ _08490_/Q _08512_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_07442_ _07446_/CLK line[113] VGND VGND VPWR VPWR _07443_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__04917__A A_h[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07373_ _07373_/A _07392_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12556__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09112_ _09116_/CLK line[123] VGND VGND VPWR VPWR _09113_/A sky130_fd_sc_hd__dfxtp_1
X_06324_ _06320_/CLK line[114] VGND VGND VPWR VPWR _06324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09043_ _09042_/Q _09072_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_06255_ _06254_/Q _06272_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09865__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05206_ _05214_/CLK line[115] VGND VGND VPWR VPWR _05206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06186_ _06186_/CLK line[51] VGND VGND VPWR VPWR _06186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05137_ _05136_/Q _05152_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10804__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VOBUF OVHB\[9\].V/Q OVHB\[9\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ _09945_/CLK _09946_/X VGND VGND VPWR VPWR _09925_/CLK sky130_fd_sc_hd__dlclkp_1
X_05068_ _05058_/CLK line[52] VGND VGND VPWR VPWR _05068_/Q sky130_fd_sc_hd__dfxtp_1
X_09876_ _09912_/A wr VGND VGND VPWR VPWR _09876_/X sky130_fd_sc_hd__and2_1
X_08827_ _13922_/X VGND VGND VPWR VPWR _08827_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08758_ _08762_/CLK line[80] VGND VGND VPWR VPWR _08759_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07709_ _07708_/Q _07742_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
X_08689_ _08688_/Q _08722_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10720_ _10728_/CLK line[90] VGND VGND VPWR VPWR _10720_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[9\].FF OVHB\[18\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[18\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10651_ _10650_/Q _10682_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11370__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06464__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13370_ _13370_/A _13377_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_10582_ _10594_/CLK line[27] VGND VGND VPWR VPWR _10583_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12321_ _12311_/CLK line[40] VGND VGND VPWR VPWR _12321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09775__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06761__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[9\].VALID\[8\].TOBUF OVHB\[9\].VALID\[8\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_12252_ _12251_/Q _12257_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13297__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11203_ _11191_/CLK line[41] VGND VGND VPWR VPWR _11204_/A sky130_fd_sc_hd__dfxtp_1
X_12183_ _12177_/CLK line[105] VGND VGND VPWR VPWR _12184_/A sky130_fd_sc_hd__dfxtp_1
X_11134_ _11133_/Q _11137_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[22\]_A0 _10883_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11065_ _11065_/CLK _11066_/X VGND VGND VPWR VPWR _11063_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_1_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10016_ _10192_/A wr VGND VGND VPWR VPWR _10016_/X sky130_fd_sc_hd__and2_1
XFILLER_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[21\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11545__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[2\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06639__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09015__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11967_ _11945_/CLK line[6] VGND VGND VPWR VPWR _11967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[2\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06936__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13706_ _13706_/A _13727_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10918_ _10918_/A _10927_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08854__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[14\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11898_ _11898_/A _11907_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_13637_ _13631_/CLK line[1] VGND VGND VPWR VPWR _13638_/A sky130_fd_sc_hd__dfxtp_1
X_10849_ _10843_/CLK line[7] VGND VGND VPWR VPWR _10850_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11280__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13568_ _13567_/Q _13587_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12519_ _12523_/CLK line[2] VGND VGND VPWR VPWR _12520_/A sky130_fd_sc_hd__dfxtp_1
X_13499_ _13497_/CLK line[66] VGND VGND VPWR VPWR _13499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06040_ _06050_/CLK line[127] VGND VGND VPWR VPWR _06040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07991_ _07990_/Q _08022_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[11\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09730_ _09730_/A _09737_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06942_ _06960_/CLK line[27] VGND VGND VPWR VPWR _06942_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[3\].TOBUF OVHB\[16\].VALID\[3\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_09661_ _09659_/CLK line[104] VGND VGND VPWR VPWR _09661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06873_ _06872_/Q _06902_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11455__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08612_ _08611_/Q _08617_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_05824_ _05836_/CLK line[28] VGND VGND VPWR VPWR _05824_/Q sky130_fd_sc_hd__dfxtp_1
X_09592_ _09592_/A _09597_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05453__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08543_ _08541_/CLK line[105] VGND VGND VPWR VPWR _08544_/A sky130_fd_sc_hd__dfxtp_1
X_05755_ _05754_/Q _05782_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13670__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08764__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08474_ _08473_/Q _08477_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05686_ _05708_/CLK line[93] VGND VGND VPWR VPWR _05687_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _07425_/CLK _07426_/X VGND VGND VPWR VPWR _07393_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12286__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07356_ _13918_/X wr VGND VGND VPWR VPWR _07356_/X sky130_fd_sc_hd__and2_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06307_ _06272_/A VGND VGND VPWR VPWR _06307_/Y sky130_fd_sc_hd__inv_2
X_07287_ _13918_/X VGND VGND VPWR VPWR _07287_/Y sky130_fd_sc_hd__inv_2
X_09026_ _09026_/A _09037_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_06238_ _06244_/CLK line[80] VGND VGND VPWR VPWR _06238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10534__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06169_ _06168_/Q _06202_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05628__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08004__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13845__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09928_ _09927_/Q _09947_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08939__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07843__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08301__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09859_ _09849_/CLK line[66] VGND VGND VPWR VPWR _09860_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12870_ _12869_/Q _12887_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05363__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11821_ _11823_/CLK line[67] VGND VGND VPWR VPWR _11821_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[27\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11752_ _11751_/Q _11767_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[18\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10707_/CLK line[68] VGND VGND VPWR VPWR _10703_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12196__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10709__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11691_/CLK line[4] VGND VGND VPWR VPWR _11684_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[2\].TOBUF OVHB\[22\].VALID\[2\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06194__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13422_ _13421_/Q _13447_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_10634_ _10634_/A _10647_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13353_ _13347_/CLK line[14] VGND VGND VPWR VPWR _13353_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[23\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10565_ _10571_/CLK line[5] VGND VGND VPWR VPWR _10565_/Q sky130_fd_sc_hd__dfxtp_1
X_12304_ _12303_/Q _12327_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13284_ _13283_/Q _13307_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_10496_ _10495_/Q _10507_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_12235_ _12227_/CLK line[15] VGND VGND VPWR VPWR _12236_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10444__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05538__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12166_ _12165_/Q _12187_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11117_ _11111_/CLK line[1] VGND VGND VPWR VPWR _11118_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12097_ _12109_/CLK line[65] VGND VGND VPWR VPWR _12098_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07753__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11048_ _11047_/Q _11067_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06369__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[13\].FF OVHB\[27\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[27\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05851__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12999_ _12999_/CLK line[108] VGND VGND VPWR VPWR _13000_/A sky130_fd_sc_hd__dfxtp_1
X_05540_ _05568_/CLK line[26] VGND VGND VPWR VPWR _05541_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10619__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05471_ _05470_/Q _05502_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_07210_ _07209_/Q _07217_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_08190_ _08189_/Q _08197_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_07141_ _07117_/CLK line[104] VGND VGND VPWR VPWR _07141_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].V OVHB\[5\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[5\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12834__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[8\].TOBUF OVHB\[14\].VALID\[8\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07928__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07072_ _07072_/A _07077_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06023_ _06023_/CLK line[105] VGND VGND VPWR VPWR _06023_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[4\].FF OVHB\[9\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[9\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07974_ _07974_/A _07987_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09713_ _09721_/CLK line[14] VGND VGND VPWR VPWR _09714_/A sky130_fd_sc_hd__dfxtp_1
X_06925_ _06923_/CLK line[5] VGND VGND VPWR VPWR _06925_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11185__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06279__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09644_ _09644_/A _09667_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06856_ _06855_/Q _06867_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05183__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[12\].TOBUF OVHB\[9\].VALID\[12\].FF/Q OVHB\[9\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05807_ _05799_/CLK line[6] VGND VGND VPWR VPWR _05807_/Q sky130_fd_sc_hd__dfxtp_1
X_09575_ _09577_/CLK line[79] VGND VGND VPWR VPWR _09575_/Q sky130_fd_sc_hd__dfxtp_1
X_06787_ _06775_/CLK line[70] VGND VGND VPWR VPWR _06788_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[4\]_A0 _10844_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08526_ _08526_/A _08547_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08494__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05738_ _05737_/Q _05747_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08473_/CLK line[65] VGND VGND VPWR VPWR _08457_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05669_ _05671_/CLK line[71] VGND VGND VPWR VPWR _05670_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07408_ _07407_/Q _07427_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08388_ _08388_/A _08407_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07339_ _07327_/CLK line[66] VGND VGND VPWR VPWR _07339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06742__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10350_ _10349_/Q _10367_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09009_ _09005_/CLK line[76] VGND VGND VPWR VPWR _09009_/Q sky130_fd_sc_hd__dfxtp_1
X_10281_ _10277_/CLK line[3] VGND VGND VPWR VPWR _10281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05358__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _12019_/Q _12047_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[2\].VALID\[11\].TOBUF OVHB\[2\].VALID\[11\].FF/Q OVHB\[2\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13575__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08669__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[20\].VALID\[7\].TOBUF OVHB\[20\].VALID\[7\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_116_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13971_ A_h[6] VGND VGND VPWR VPWR _13979_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[7\].VALID\[6\].FF OVHB\[7\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[7\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08966__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12922_ _12992_/A VGND VGND VPWR VPWR _12922_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[18\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05093__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12853_ _12881_/CLK line[32] VGND VGND VPWR VPWR _12853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11823__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11804_ _11803_/Q _11837_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06917__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12784_ _12783_/Q _12817_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _11757_/CLK line[42] VGND VGND VPWR VPWR _11735_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11665_/Q _11697_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13405_/A _13412_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_10617_ _10627_/CLK line[43] VGND VGND VPWR VPWR _10617_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _11605_/CLK line[107] VGND VGND VPWR VPWR _11597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[18\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13336_ _13308_/CLK line[120] VGND VGND VPWR VPWR _13336_/Q sky130_fd_sc_hd__dfxtp_1
X_10548_ _10547_/Q _10577_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10174__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13267_ _13266_/Q _13272_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_10479_ _10473_/CLK line[108] VGND VGND VPWR VPWR _10479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10752__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05268__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12218_ _12204_/CLK line[121] VGND VGND VPWR VPWR _12218_/Q sky130_fd_sc_hd__dfxtp_1
X_13198_ _13194_/CLK line[57] VGND VGND VPWR VPWR _13198_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[21\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10471__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13485__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12149_ _12148_/Q _12152_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07483__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04971_ _04947_/CLK line[8] VGND VGND VPWR VPWR _04971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06710_ _06709_/Q _06727_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07690_ _07689_/Q _07707_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].V OVHB\[10\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[10\].V/Q sky130_fd_sc_hd__dfrtp_1
X_06641_ _06633_/CLK line[3] VGND VGND VPWR VPWR _06641_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11733__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09360_ _09360_/A _09387_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_06572_ _06571_/Q _06587_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05731__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08311_ _08329_/CLK line[13] VGND VGND VPWR VPWR _08311_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[8\].FF OVHB\[5\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[5\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10349__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05523_ _05519_/CLK line[4] VGND VGND VPWR VPWR _05524_/A sky130_fd_sc_hd__dfxtp_1
X_09291_ _09307_/CLK line[77] VGND VGND VPWR VPWR _09291_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10927__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ _08241_/Q _08267_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_05454_ _05453_/Q _05467_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10646__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12564__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05385_ _05391_/CLK line[69] VGND VGND VPWR VPWR _05385_/Q sky130_fd_sc_hd__dfxtp_1
X_08173_ _08175_/CLK line[78] VGND VGND VPWR VPWR _08173_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[2\].TOBUF OVHB\[29\].VALID\[2\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07658__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07124_ _07123_/Q _07147_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07055_ _07043_/CLK line[79] VGND VGND VPWR VPWR _07056_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09873__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06006_ _06006_/A _06027_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[23\].VALID\[11\].FF OVHB\[23\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[23\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11908__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10812__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07393__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05906__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07957_ _07981_/CLK line[107] VGND VGND VPWR VPWR _07958_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[25\].VALID\[13\].TOBUF OVHB\[25\].VALID\[13\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_06908_ _06907_/Q _06937_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06587__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07888_ _07887_/Q _07917_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09627_ _09626_/Q _09632_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12739__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06839_ _06839_/CLK line[108] VGND VGND VPWR VPWR _06839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09558_ _09554_/CLK line[57] VGND VGND VPWR VPWR _09558_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08509_ _08508_/Q _08512_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09489_ _09489_/A _09492_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11520_ _11520_/CLK _11521_/X VGND VGND VPWR VPWR _11500_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _11592_/A wr VGND VGND VPWR VPWR _11451_/X sky130_fd_sc_hd__and2_1
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[13\].FF OVHB\[13\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[13\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07568__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06472__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10402_ _13931_/X VGND VGND VPWR VPWR _10402_/Y sky130_fd_sc_hd__inv_2
X_11382_ _11311_/A VGND VGND VPWR VPWR _11382_/Y sky130_fd_sc_hd__inv_2
X_13121_ _13121_/A _13132_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_10333_ _10341_/CLK line[32] VGND VGND VPWR VPWR _10333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09783__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13052_ _13050_/CLK line[118] VGND VGND VPWR VPWR _13052_/Q sky130_fd_sc_hd__dfxtp_1
X_10264_ _10263_/Q _10297_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12003_ _12003_/A _12012_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10722__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10195_ _10217_/CLK line[106] VGND VGND VPWR VPWR _10195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08399__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07881__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _13950_/A _13950_/B _13950_/C _13957_/D VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__and4bb_4
X_12905_ _12904_/Q _12922_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12649__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13885_ _13884_/Q _13902_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11553__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12011__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06647__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12836_ _12820_/CLK line[19] VGND VGND VPWR VPWR _12836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09023__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12767_ _12766_/Q _12782_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09958__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11718_ _11706_/CLK line[20] VGND VGND VPWR VPWR _11719_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[0\].FF OVHB\[14\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[14\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12698_ _12708_/CLK line[84] VGND VGND VPWR VPWR _12698_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[4\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11649_ _11649_/A _11662_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[4\].FF OVHB\[31\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[31\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05170_ _05170_/A _05187_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06382__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13319_ _13318_/Q _13342_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11728__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08860_ _08860_/CLK _08861_/X VGND VGND VPWR VPWR _08850_/CLK sky130_fd_sc_hd__dlclkp_1
X_07811_ _13920_/X wr VGND VGND VPWR VPWR _07811_/X sky130_fd_sc_hd__and2_1
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08791_ _13922_/X wr VGND VGND VPWR VPWR _08791_/X sky130_fd_sc_hd__and2_1
XOVHB\[2\].VALID\[4\].TOBUF OVHB\[2\].VALID\[4\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_07742_ _07672_/A VGND VGND VPWR VPWR _07742_/Y sky130_fd_sc_hd__inv_2
X_04954_ _04953_/Q _04977_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[7\].TOBUF OVHB\[27\].VALID\[7\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07673_ _07679_/CLK line[96] VGND VGND VPWR VPWR _07673_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11463__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09412_ _09414_/CLK line[118] VGND VGND VPWR VPWR _09412_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06557__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06624_ _06623_/Q _06657_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05461__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10079__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09343_ _09343_/A _09352_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_06555_ _06565_/CLK line[106] VGND VGND VPWR VPWR _06556_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[1\]_A3 _13568_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05506_ _05505_/Q _05537_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08772__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09274_ _09256_/CLK line[55] VGND VGND VPWR VPWR _09274_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08127__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06486_ _06485_/Q _06517_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08225_ _08224_/Q _08232_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_05437_ _05445_/CLK line[107] VGND VGND VPWR VPWR _05438_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].CGAND _13909_/X wr VGND VGND VPWR VPWR OVHB\[11\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__07388__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08156_ _08134_/CLK line[56] VGND VGND VPWR VPWR _08156_/Q sky130_fd_sc_hd__dfxtp_1
X_05368_ _05367_/Q _05397_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_07107_ _07106_/Q _07112_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_05299_ _05299_/CLK line[44] VGND VGND VPWR VPWR _05300_/A sky130_fd_sc_hd__dfxtp_1
X_08087_ _08086_/Q _08092_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[2\].FF OVHB\[12\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[12\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07038_ _07030_/CLK line[57] VGND VGND VPWR VPWR _07038_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11638__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05636__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09108__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08012__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08989_ _08988_/Q _09002_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13853__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08947__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10951_ _10950_/Q _10962_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13670_ _13682_/CLK line[31] VGND VGND VPWR VPWR _13670_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05371__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10882_ _10872_/CLK line[22] VGND VGND VPWR VPWR _10882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ _12621_/A _12642_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09421__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _12560_/CLK line[17] VGND VGND VPWR VPWR _12552_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11502_/Q _11522_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12482_/Q _12502_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12782__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07298__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ _11440_/CLK line[18] VGND VGND VPWR VPWR _11434_/Q sky130_fd_sc_hd__dfxtp_1
X_11365_ _11364_/Q _11382_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05396__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13104_ _13120_/CLK line[28] VGND VGND VPWR VPWR _13104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10316_ _10314_/CLK line[19] VGND VGND VPWR VPWR _10316_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[7\].FF OVHB\[28\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[28\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11296_ _11302_/CLK line[83] VGND VGND VPWR VPWR _11297_/A sky130_fd_sc_hd__dfxtp_1
X_13035_ _13034_/Q _13062_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10452__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10247_ _10246_/Q _10262_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05546__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10178_ _10188_/CLK line[84] VGND VGND VPWR VPWR _10178_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13763__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[4\].FF OVHB\[10\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[10\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07761__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12379__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13937_ A[5] VGND VGND VPWR VPWR _13946_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12957__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13868_ _13882_/CLK line[112] VGND VGND VPWR VPWR _13868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12676__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _12819_/A _12852_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_13799_ _13798_/Q _13832_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09688__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06340_ _06340_/CLK _06341_/X VGND VGND VPWR VPWR _06320_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_72_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10627__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06271_ _06272_/A wr VGND VGND VPWR VPWR _06271_/X sky130_fd_sc_hd__and2_1
XDATA\[29\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _10925_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13003__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[9\].TOBUF OVHB\[0\].VALID\[9\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_08010_ _08000_/CLK line[117] VGND VGND VPWR VPWR _08010_/Q sky130_fd_sc_hd__dfxtp_1
X_05222_ _05152_/A VGND VGND VPWR VPWR _05222_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07001__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05153_ _05157_/CLK line[96] VGND VGND VPWR VPWR _05153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12842__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11101__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07936__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09961_ _09960_/Q _09982_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_05084_ _05083_/Q _05117_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_08912_ _08922_/CLK line[17] VGND VGND VPWR VPWR _08912_/Q sky130_fd_sc_hd__dfxtp_1
X_09892_ _09908_/CLK line[81] VGND VGND VPWR VPWR _09892_/Q sky130_fd_sc_hd__dfxtp_1
X_08843_ _08843_/A _08862_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_08774_ _08762_/CLK line[82] VGND VGND VPWR VPWR _08775_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05986_ _05984_/CLK line[88] VGND VGND VPWR VPWR _05986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[26\].VALID\[9\].FF OVHB\[26\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[26\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07725_ _07725_/A _07742_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_04937_ A_h[14] _04937_/B2 A_h[14] _04937_/B2 VGND VGND VPWR VPWR _04937_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11193__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06287__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07656_ _07644_/CLK line[83] VGND VGND VPWR VPWR _07656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[5\].VOBUF OVHB\[5\].V/Q OVHB\[5\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06607_ _06606_/Q _06622_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_07587_ _07587_/A _07602_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09598__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09326_ _09320_/CLK line[93] VGND VGND VPWR VPWR _09327_/A sky130_fd_sc_hd__dfxtp_1
X_06538_ _06528_/CLK line[84] VGND VGND VPWR VPWR _06538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09257_ _09257_/A _09282_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_06469_ _06468_/Q _06482_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_08208_ _08208_/CLK line[94] VGND VGND VPWR VPWR _08209_/A sky130_fd_sc_hd__dfxtp_1
X_09188_ _09200_/CLK line[30] VGND VGND VPWR VPWR _09188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[17\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08139_ _08138_/Q _08162_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12752__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06750__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11150_ _11148_/CLK line[31] VGND VGND VPWR VPWR _11150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11368__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10101_ _10100_/Q _10122_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_11081_ _11080_/Q _11102_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[18\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _07670_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_89_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[15\].VALID\[11\].TOBUF OVHB\[15\].VALID\[11\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10032_ _10042_/CLK line[17] VGND VGND VPWR VPWR _10032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13583__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08677__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11983_ _11982_/Q _12012_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[9\].VALID\[4\].TOBUF OVHB\[9\].VALID\[4\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_1_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13722_ _13721_/Q _13727_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10934_ _10930_/CLK line[60] VGND VGND VPWR VPWR _10934_/Q sky130_fd_sc_hd__dfxtp_1
X_13653_ _13631_/CLK line[9] VGND VGND VPWR VPWR _13653_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12927__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10297__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10865_ _10864_/Q _10892_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11831__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12604_ _12603_/Q _12607_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06925__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[13\].FF OVHB\[4\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[4\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13584_ _13584_/A _13587_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10796_ _10804_/CLK line[125] VGND VGND VPWR VPWR _10796_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09301__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12535_ _12535_/CLK _12536_/X VGND VGND VPWR VPWR _12523_/CLK sky130_fd_sc_hd__dlclkp_1
X_12466_ _13943_/X wr VGND VGND VPWR VPWR _12466_/X sky130_fd_sc_hd__and2_1
XFILLER_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13758__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11417_ _11592_/A VGND VGND VPWR VPWR _11417_/Y sky130_fd_sc_hd__inv_2
X_12397_ _13943_/X VGND VGND VPWR VPWR _12397_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06660__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11348_ _11370_/CLK line[112] VGND VGND VPWR VPWR _11348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11278__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10182__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11279_ _11278_/Q _11312_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05276__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13018_ _13017_/Q _13027_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13493__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08587__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05840_ _05836_/CLK line[21] VGND VGND VPWR VPWR _05841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07491__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _07285_/CLK sky130_fd_sc_hd__clkbuf_4
X_05771_ _05771_/A _05782_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_07510_ _07518_/CLK line[31] VGND VGND VPWR VPWR _07510_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11591__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08490_ _08480_/CLK line[95] VGND VGND VPWR VPWR _08490_/Q sky130_fd_sc_hd__dfxtp_1
X_07441_ _07440_/Q _07462_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11741__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06835__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07372_ _07380_/CLK line[81] VGND VGND VPWR VPWR _07373_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09111_ _09111_/A _09142_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10357__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06323_ _06322_/Q _06342_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_09042_ _09068_/CLK line[91] VGND VGND VPWR VPWR _09042_/Q sky130_fd_sc_hd__dfxtp_1
X_06254_ _06244_/CLK line[82] VGND VGND VPWR VPWR _06254_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[11\].FF OVHB\[28\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[28\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13668__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05205_ _05204_/Q _05222_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_06185_ _06184_/Q _06202_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07666__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05136_ _05122_/CLK line[83] VGND VGND VPWR VPWR _05136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10092__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11766__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09944_ _09944_/A _09947_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_05067_ _05066_/Q _05082_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09875_ _09875_/CLK _09876_/X VGND VGND VPWR VPWR _09849_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11916__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13981__A A_h[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08826_ _13922_/X wr VGND VGND VPWR VPWR _08826_/X sky130_fd_sc_hd__and2_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05914__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08757_ _13922_/X VGND VGND VPWR VPWR _08757_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05969_ _05968_/Q _05992_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_07708_ _07724_/CLK line[112] VGND VGND VPWR VPWR _07708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08688_ _08710_/CLK line[48] VGND VGND VPWR VPWR _08688_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[31\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[13\].FF OVHB\[18\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[18\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07639_ _07638_/Q _07672_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_10650_ _10656_/CLK line[58] VGND VGND VPWR VPWR _10650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09309_ _09307_/CLK line[71] VGND VGND VPWR VPWR _09309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10267__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10581_ _10580_/Q _10612_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12320_ _12320_/A _12327_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12251_ _12227_/CLK line[8] VGND VGND VPWR VPWR _12251_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12482__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07576__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[9\].TOBUF OVHB\[7\].VALID\[9\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_11202_ _11202_/A _11207_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12182_ _12182_/A _12187_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11098__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11133_ _11111_/CLK line[9] VGND VGND VPWR VPWR _11133_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09791__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[22\]_A1 _13473_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11064_ _11064_/A _11067_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10015_ _10015_/CLK _10016_/X VGND VGND VPWR VPWR _10011_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10730__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05824__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08200__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DEC.DEC0.AND3_A A[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11966_ _11965_/Q _11977_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_13705_ _13701_/CLK line[47] VGND VGND VPWR VPWR _13706_/A sky130_fd_sc_hd__dfxtp_1
X_10917_ _10903_/CLK line[38] VGND VGND VPWR VPWR _10918_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12657__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11897_ _11901_/CLK line[102] VGND VGND VPWR VPWR _11898_/A sky130_fd_sc_hd__dfxtp_1
X_13636_ _13635_/Q _13657_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[7\] _11410_/Z _05600_/Z _13510_/Z _07140_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[7] sky130_fd_sc_hd__mux4_1
X_10848_ _10848_/A _10857_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09031__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13567_ _13559_/CLK line[97] VGND VGND VPWR VPWR _13567_/Q sky130_fd_sc_hd__dfxtp_1
X_10779_ _10783_/CLK line[103] VGND VGND VPWR VPWR _10779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09966__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13131__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12518_ _12517_/Q _12537_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_13498_ _13498_/A _13517_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12449_ _12449_/CLK line[98] VGND VGND VPWR VPWR _12449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10905__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06390__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07990_ _08000_/CLK line[122] VGND VGND VPWR VPWR _07990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06941_ _06940_/Q _06972_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09660_ _09660_/A _09667_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_06872_ _06892_/CLK line[123] VGND VGND VPWR VPWR _06872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09206__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[4\].TOBUF OVHB\[14\].VALID\[4\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_08611_ _08609_/CLK line[8] VGND VGND VPWR VPWR _08611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[0\].VALID\[11\].FF OVHB\[0\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[0\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05823_ _05822_/Q _05852_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09591_ _09577_/CLK line[72] VGND VGND VPWR VPWR _09592_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08542_ _08542_/A _08547_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13306__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05754_ _05756_/CLK line[124] VGND VGND VPWR VPWR _05754_/Q sky130_fd_sc_hd__dfxtp_1
X_08473_ _08473_/CLK line[73] VGND VGND VPWR VPWR _08473_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11471__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05685_ _05685_/A _05712_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07424_ _07423_/Q _07427_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06565__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07355_ _07355_/CLK _07356_/X VGND VGND VPWR VPWR _07327_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_137_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06306_ _06272_/A wr VGND VGND VPWR VPWR _06306_/X sky130_fd_sc_hd__and2_1
XANTENNA__08780__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07286_ _13918_/X wr VGND VGND VPWR VPWR _07286_/X sky130_fd_sc_hd__and2_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13398__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09025_ _09005_/CLK line[69] VGND VGND VPWR VPWR _09026_/A sky130_fd_sc_hd__dfxtp_1
X_06237_ _06272_/A VGND VGND VPWR VPWR _06237_/Y sky130_fd_sc_hd__inv_2
X_06168_ _06186_/CLK line[48] VGND VGND VPWR VPWR _06168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[10\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05119_ _05118_/Q _05152_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_06099_ _06098_/Q _06132_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_09927_ _09925_/CLK line[97] VGND VGND VPWR VPWR _09927_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11646__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09858_ _09857_/Q _09877_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[17\].CG clk OVHB\[17\].CGAND/X VGND VGND VPWR VPWR OVHB\[17\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_85_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[9\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09116__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08809_ _08823_/CLK line[98] VGND VGND VPWR VPWR _08809_/Q sky130_fd_sc_hd__dfxtp_1
X_09789_ _09793_/CLK line[34] VGND VGND VPWR VPWR _09789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13861__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _11820_/A _11837_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08955__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11751_ _11757_/CLK line[35] VGND VGND VPWR VPWR _11751_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10702_/A _10717_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[3\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11682_ _11681_/Q _11697_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13439_/CLK line[45] VGND VGND VPWR VPWR _13421_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10627_/CLK line[36] VGND VGND VPWR VPWR _10634_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[3\].TOBUF OVHB\[20\].VALID\[3\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08690__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13352_ _13351_/Q _13377_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_10564_ _10564_/A _10577_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_12303_ _12311_/CLK line[46] VGND VGND VPWR VPWR _12303_/Q sky130_fd_sc_hd__dfxtp_1
X_13283_ _13285_/CLK line[110] VGND VGND VPWR VPWR _13283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10495_ _10473_/CLK line[101] VGND VGND VPWR VPWR _10495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12234_ _12233_/Q _12257_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12165_ _12177_/CLK line[111] VGND VGND VPWR VPWR _12165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11116_ _11116_/A _11137_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12096_ _12095_/Q _12117_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[11\].FF OVHB\[14\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[14\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10460__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11047_ _11063_/CLK line[97] VGND VGND VPWR VPWR _11047_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05554__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13771__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08865__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05851__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _12997_/Q _13027_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12387__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11949_ _11945_/CLK line[12] VGND VGND VPWR VPWR _11949_/Q sky130_fd_sc_hd__dfxtp_1
X_05470_ _05476_/CLK line[122] VGND VGND VPWR VPWR _05470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13619_ _13618_/Q _13622_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09696__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07140_ _07139_/Q _07147_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[11\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13796__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10635__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07071_ _07043_/CLK line[72] VGND VGND VPWR VPWR _07072_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[9\].TOBUF OVHB\[12\].VALID\[9\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13011__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05729__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06022_ _06022_/A _06027_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08105__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[13\].TOBUF OVHB\[5\].VALID\[13\].FF/Q OVHB\[5\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07944__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07973_ _07981_/CLK line[100] VGND VGND VPWR VPWR _07974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10370__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09712_ _09711_/Q _09737_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[8\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _13585_/CLK sky130_fd_sc_hd__clkbuf_4
X_06924_ _06923_/Q _06937_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_09643_ _09659_/CLK line[110] VGND VGND VPWR VPWR _09644_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06855_ _06839_/CLK line[101] VGND VGND VPWR VPWR _06855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05806_ _05805_/Q _05817_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09574_ _09573_/Q _09597_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_06786_ _06785_/Q _06797_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[4\]_A1 _05594_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08525_ _08541_/CLK line[111] VGND VGND VPWR VPWR _08526_/A sky130_fd_sc_hd__dfxtp_1
X_05737_ _05739_/CLK line[102] VGND VGND VPWR VPWR _05737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12297__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06295__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _08456_/A _08477_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_05668_ _05668_/A _05677_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _07393_/CLK line[97] VGND VGND VPWR VPWR _07407_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[12\]_A0 _10830_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _08383_/CLK line[33] VGND VGND VPWR VPWR _08388_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05599_ _05575_/CLK line[39] VGND VGND VPWR VPWR _05599_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[28\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07338_ _07337_/Q _07357_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10545__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07269_ _07267_/CLK line[34] VGND VGND VPWR VPWR _07269_/Q sky130_fd_sc_hd__dfxtp_1
X_09008_ _09007_/Q _09037_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_10280_ _10279_/Q _10297_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12760__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07854__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11376__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ A_h[5] VGND VGND VPWR VPWR _13979_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12921_ _12992_/A wr VGND VGND VPWR VPWR _12921_/X sky130_fd_sc_hd__and2_1
XFILLER_24_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[9\].VALID\[13\].FF OVHB\[9\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[9\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[31\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12852_ _12992_/A VGND VGND VPWR VPWR _12852_/Y sky130_fd_sc_hd__inv_2
XOVHB\[22\].VALID\[0\].FF OVHB\[22\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[22\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _13200_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11803_ _11823_/CLK line[64] VGND VGND VPWR VPWR _11803_/Q sky130_fd_sc_hd__dfxtp_1
X_12783_ _12803_/CLK line[0] VGND VGND VPWR VPWR _12783_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12000__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11734_ _11733_/Q _11767_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11691_/CLK line[10] VGND VGND VPWR VPWR _11665_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12935__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[24\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ _10615_/Q _10647_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06933__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13404_ _13394_/CLK line[23] VGND VGND VPWR VPWR _13405_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _11595_/Q _11627_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13334_/Q _13342_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_10547_ _10571_/CLK line[11] VGND VGND VPWR VPWR _10547_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ _13254_/CLK line[88] VGND VGND VPWR VPWR _13266_/Q sky130_fd_sc_hd__dfxtp_1
X_10478_ _10477_/Q _10507_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_12217_ _12216_/Q _12222_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_13197_ _13197_/A _13202_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12148_ _12130_/CLK line[89] VGND VGND VPWR VPWR _12148_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11286__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[27\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _10540_/CLK sky130_fd_sc_hd__clkbuf_4
X_12079_ _12078_/Q _12082_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_04970_ _04969_/Q _04977_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05284__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08595__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06640_ _06639_/Q _06657_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06571_ _06565_/CLK line[99] VGND VGND VPWR VPWR _06571_/Q sky130_fd_sc_hd__dfxtp_1
X_08310_ _08309_/Q _08337_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_05522_ _05521_/Q _05537_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09290_ _09289_/Q _09317_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08241_ _08257_/CLK line[109] VGND VGND VPWR VPWR _08241_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[6\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _12815_/CLK sky130_fd_sc_hd__clkbuf_4
X_05453_ _05445_/CLK line[100] VGND VGND VPWR VPWR _05453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[20\].VALID\[2\].FF OVHB\[20\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[20\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[0\].TOBUF OVHB\[2\].VALID\[0\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06843__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _08172_/A _08197_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05384_ _05384_/A _05397_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_07123_ _07117_/CLK line[110] VGND VGND VPWR VPWR _07123_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[3\].TOBUF OVHB\[27\].VALID\[3\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_118_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05459__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07054_ _07053_/Q _07077_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[14\].TOBUF OVHB\[21\].VALID\[14\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_86_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13676__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06005_ _06023_/CLK line[111] VGND VGND VPWR VPWR _06006_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[17\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[5\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07956_ _07956_/A _07987_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05194__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06907_ _06923_/CLK line[11] VGND VGND VPWR VPWR _06907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07887_ _07905_/CLK line[75] VGND VGND VPWR VPWR _07887_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11924__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09626_ _09626_/CLK line[88] VGND VGND VPWR VPWR _09626_/Q sky130_fd_sc_hd__dfxtp_1
X_06838_ _06837_/Q _06867_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _10155_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09557_ _09557_/A _09562_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_06769_ _06775_/CLK line[76] VGND VGND VPWR VPWR _06770_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08508_ _08480_/CLK line[89] VGND VGND VPWR VPWR _08508_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09488_ _09482_/CLK line[25] VGND VGND VPWR VPWR _09489_/A sky130_fd_sc_hd__dfxtp_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[19\].VALID\[3\].FF OVHB\[19\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[19\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _08438_/Q _08442_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[25\] _10329_/Z _07039_/Z _13549_/Z _07179_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[25] sky130_fd_sc_hd__mux4_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11450_ _11450_/CLK _11451_/X VGND VGND VPWR VPWR _11440_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _13931_/X wr VGND VGND VPWR VPWR _10401_/X sky130_fd_sc_hd__and2_1
XANTENNA__05012__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10275__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11381_ _11311_/A wr VGND VGND VPWR VPWR _11381_/X sky130_fd_sc_hd__and2_1
XANTENNA__05369__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _13120_/CLK line[21] VGND VGND VPWR VPWR _13121_/A sky130_fd_sc_hd__dfxtp_1
X_10332_ _13931_/X VGND VGND VPWR VPWR _10332_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[26\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12490__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13051_ _13050_/Q _13062_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10263_ _10277_/CLK line[0] VGND VGND VPWR VPWR _10263_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[9\].TOBUF OVHB\[19\].VALID\[9\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07584__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12002_ _12002_/CLK line[22] VGND VGND VPWR VPWR _12003_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10194_ _10193_/Q _10227_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07881__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13953_ _13950_/C _13950_/B _13950_/A _13957_/D VGND VGND VPWR VPWR _13953_/X sky130_fd_sc_hd__and4b_4
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12904_ _12902_/CLK line[50] VGND VGND VPWR VPWR _12904_/Q sky130_fd_sc_hd__dfxtp_1
X_13884_ _13882_/CLK line[114] VGND VGND VPWR VPWR _13884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05832__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12835_ _12835_/A _12852_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12774_/CLK line[115] VGND VGND VPWR VPWR _12766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[25\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _09770_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12665__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11717_ _11716_/Q _11732_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12697_ _12696_/Q _12712_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07759__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _11636_/CLK line[116] VGND VGND VPWR VPWR _11649_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[15\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _06900_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_11_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11579_ _11578_/Q _11592_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09974__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13318_ _13308_/CLK line[126] VGND VGND VPWR VPWR _13318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[17\].VALID\[5\].FF OVHB\[17\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[17\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10913__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13249_ _13248_/Q _13272_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[5\].VALID\[11\].FF OVHB\[5\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[5\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07810_ _07810_/CLK _07811_/X VGND VGND VPWR VPWR _07788_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08790_ _08790_/CLK _08791_/X VGND VGND VPWR VPWR _08762_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_38_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07741_ _07672_/A wr VGND VGND VPWR VPWR _07741_/X sky130_fd_sc_hd__and2_1
XOVHB\[0\].VALID\[5\].TOBUF OVHB\[0\].VALID\[5\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_04953_ _04947_/CLK line[14] VGND VGND VPWR VPWR _04953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07672_ _07672_/A VGND VGND VPWR VPWR _07672_/Y sky130_fd_sc_hd__inv_2
XOVHB\[25\].VALID\[8\].TOBUF OVHB\[25\].VALID\[8\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09411_ _09410_/Q _09422_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_06623_ _06633_/CLK line[0] VGND VGND VPWR VPWR _06623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09342_ _09320_/CLK line[86] VGND VGND VPWR VPWR _09343_/A sky130_fd_sc_hd__dfxtp_1
X_06554_ _06553_/Q _06587_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_05505_ _05519_/CLK line[10] VGND VGND VPWR VPWR _05505_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12575__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09273_ _09272_/Q _09282_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_06485_ _06489_/CLK line[74] VGND VGND VPWR VPWR _06485_/Q sky130_fd_sc_hd__dfxtp_1
X_08224_ _08208_/CLK line[87] VGND VGND VPWR VPWR _08224_/Q sky130_fd_sc_hd__dfxtp_1
X_05436_ _05436_/A _05467_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06573__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08155_ _08154_/Q _08162_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_05367_ _05391_/CLK line[75] VGND VGND VPWR VPWR _05367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09884__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07106_ _07098_/CLK line[88] VGND VGND VPWR VPWR _07106_/Q sky130_fd_sc_hd__dfxtp_1
X_08086_ _08070_/CLK line[24] VGND VGND VPWR VPWR _08086_/Q sky130_fd_sc_hd__dfxtp_1
X_05298_ _05297_/Q _05327_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[14\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _06515_/CLK sky130_fd_sc_hd__clkbuf_4
X_07037_ _07036_/Q _07042_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10823__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[1\].VOBUF OVHB\[1\].V/Q OVHB\[1\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08988_ _08972_/CLK line[52] VGND VGND VPWR VPWR _08988_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[7\].FF OVHB\[15\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[15\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07939_ _07938_/Q _07952_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11654__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _10930_/CLK line[53] VGND VGND VPWR VPWR _10950_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06748__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09124__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09609_ _09608_/Q _09632_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09702__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10881_ _10880_/Q _10892_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08963__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12620_ _12638_/CLK line[63] VGND VGND VPWR VPWR _12621_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09421__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _12550_/Q _12572_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _11500_/CLK line[49] VGND VGND VPWR VPWR _11502_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06483__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12490_/CLK line[113] VGND VGND VPWR VPWR _12482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[7\].TOBUF OVHB\[31\].VALID\[7\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ _11432_/Q _11452_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05099__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05677__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[0\].TOBUF OVHB\[9\].VALID\[0\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[29\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11364_ _11370_/CLK line[114] VGND VGND VPWR VPWR _11364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[19\].VALID\[11\].FF OVHB\[19\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[19\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11829__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _13103_/A _13132_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_10315_ _10314_/Q _10332_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05396__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11295_ _11294_/Q _11312_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13034_ _13050_/CLK line[124] VGND VGND VPWR VPWR _13034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10246_ _10248_/CLK line[115] VGND VGND VPWR VPWR _10246_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[13\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _06130_/CLK sky130_fd_sc_hd__clkbuf_4
X_10177_ _10177_/A _10192_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11564__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06658__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13936_ A[4] VGND VGND VPWR VPWR _13944_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__05562__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867_ _13907_/X VGND VGND VPWR VPWR _13867_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08873__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12818_ _12820_/CLK line[16] VGND VGND VPWR VPWR _12819_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[9\].FF OVHB\[13\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[13\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13798_ _13822_/CLK line[80] VGND VGND VPWR VPWR _13798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12749_ _12748_/Q _12782_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07489__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06270_ _06270_/CLK _06271_/X VGND VGND VPWR VPWR _06244_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06971__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05221_ _05152_/A wr VGND VGND VPWR VPWR _05221_/X sky130_fd_sc_hd__and2_1
XFILLER_128_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05152_ _05152_/A VGND VGND VPWR VPWR _05152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11739__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10643__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11101__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09960_ _09978_/CLK line[127] VGND VGND VPWR VPWR _09960_/Q sky130_fd_sc_hd__dfxtp_1
X_05083_ _05093_/CLK line[64] VGND VGND VPWR VPWR _05083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05737__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08113__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08911_ _08910_/Q _08932_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09891_ _09890_/Q _09912_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[18\].VALID\[13\].TOBUF OVHB\[18\].VALID\[13\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_08842_ _08850_/CLK line[113] VGND VGND VPWR VPWR _08843_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08773_ _08772_/Q _08792_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_05985_ _05984_/Q _05992_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07724_ _07724_/CLK line[114] VGND VGND VPWR VPWR _07725_/A sky130_fd_sc_hd__dfxtp_1
X_04936_ _04932_/X _04936_/B _04936_/C _04935_/X VGND VGND VPWR VPWR _04942_/C sky130_fd_sc_hd__and4_4
XANTENNA__05472__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07655_ _07654_/Q _07672_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06606_ _06596_/CLK line[115] VGND VGND VPWR VPWR _06606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ _07572_/CLK line[51] VGND VGND VPWR VPWR _07587_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07042__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09325_ _09324_/Q _09352_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_06537_ _06536_/Q _06552_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10818__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07399__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09256_ _09256_/CLK line[61] VGND VGND VPWR VPWR _09257_/A sky130_fd_sc_hd__dfxtp_1
X_06468_ _06464_/CLK line[52] VGND VGND VPWR VPWR _06468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08207_ _08206_/Q _08232_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_05419_ _05418_/Q _05432_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_09187_ _09187_/A _09212_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_06399_ _06399_/A _06412_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[12\].TOBUF OVHB\[11\].VALID\[12\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_08138_ _08134_/CLK line[62] VGND VGND VPWR VPWR _08138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10553__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08069_ _08068_/Q _08092_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05647__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10100_ _10100_/CLK line[63] VGND VGND VPWR VPWR _10100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[8\].CGAND _13552_/A wr VGND VGND VPWR VPWR OVHB\[8\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__08023__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11080_ _11090_/CLK line[127] VGND VGND VPWR VPWR _11080_/Q sky130_fd_sc_hd__dfxtp_1
X_10031_ _10030_/Q _10052_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07862__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].CGAND_A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07217__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[8\].VALID\[0\].FF OVHB\[8\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[8\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06478__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11982_ _12002_/CLK line[27] VGND VGND VPWR VPWR _11982_/Q sky130_fd_sc_hd__dfxtp_1
X_13721_ _13701_/CLK line[40] VGND VGND VPWR VPWR _13721_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[5\].TOBUF OVHB\[7\].VALID\[5\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
X_10933_ _10932_/Q _10962_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09789__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13652_ _13651_/Q _13657_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_10864_ _10872_/CLK line[28] VGND VGND VPWR VPWR _10864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12603_ _12601_/CLK line[41] VGND VGND VPWR VPWR _12603_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10728__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _13559_/CLK line[105] VGND VGND VPWR VPWR _13584_/A sky130_fd_sc_hd__dfxtp_1
X_10795_ _10794_/Q _10822_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13104__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12534_ _12534_/A _12537_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07102__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12943__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12465_ _12465_/CLK _12466_/X VGND VGND VPWR VPWR _12449_/CLK sky130_fd_sc_hd__dlclkp_1
X_11416_ _11592_/A wr VGND VGND VPWR VPWR _11416_/X sky130_fd_sc_hd__and2_1
X_12396_ _13943_/X wr VGND VGND VPWR VPWR _12396_/X sky130_fd_sc_hd__and2_1
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11347_ _11311_/A VGND VGND VPWR VPWR _11347_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09029__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11278_ _11302_/CLK line[80] VGND VGND VPWR VPWR _11278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08511__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13017_ _12999_/CLK line[102] VGND VGND VPWR VPWR _13017_/Q sky130_fd_sc_hd__dfxtp_1
X_10229_ _10228_/Q _10262_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11294__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11872__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06388__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05770_ _05756_/CLK line[117] VGND VGND VPWR VPWR _05771_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11591__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13919_ _13923_/C _13922_/B _13923_/B _13923_/D VGND VGND VPWR VPWR _07672_/A sky130_fd_sc_hd__and4bb_4
XFILLER_39_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07440_ _07446_/CLK line[127] VGND VGND VPWR VPWR _07440_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[12\].TOBUF OVHB\[31\].VALID\[12\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_07371_ _07370_/Q _07392_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[2\].FF OVHB\[6\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[6\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09110_ _09116_/CLK line[122] VGND VGND VPWR VPWR _09111_/A sky130_fd_sc_hd__dfxtp_1
X_06322_ _06320_/CLK line[113] VGND VGND VPWR VPWR _06322_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07012__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09041_ _09041_/A _09072_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12853__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06253_ _06252_/Q _06272_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[0\].TOBUF OVHB\[14\].VALID\[0\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_102_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05204_ _05214_/CLK line[114] VGND VGND VPWR VPWR _05204_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06851__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06184_ _06186_/CLK line[50] VGND VGND VPWR VPWR _06184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11469__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05135_ _05135_/A _05152_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09943_ _09925_/CLK line[105] VGND VGND VPWR VPWR _09944_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11766__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05066_ _05058_/CLK line[51] VGND VGND VPWR VPWR _05066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13684__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08778__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09874_ _09873_/Q _09877_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[29\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08825_ _08825_/CLK _08826_/X VGND VGND VPWR VPWR _08823_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_39_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08756_ _13922_/X wr VGND VGND VPWR VPWR _08756_/X sky130_fd_sc_hd__and2_1
X_05968_ _05984_/CLK line[94] VGND VGND VPWR VPWR _05968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04919_ A_h[20] _04919_/B2 A_h[20] _04919_/B2 VGND VGND VPWR VPWR _04921_/C sky130_fd_sc_hd__a2bb2o_4
X_07707_ _07672_/A VGND VGND VPWR VPWR _07707_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08687_ _13922_/X VGND VGND VPWR VPWR _08687_/Y sky130_fd_sc_hd__inv_2
X_05899_ _05898_/Q _05922_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11932__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07638_ _07644_/CLK line[80] VGND VGND VPWR VPWR _07638_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09402__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07569_ _07568_/Q _07602_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_09308_ _09307_/Q _09317_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08018__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10580_ _10594_/CLK line[26] VGND VGND VPWR VPWR _10580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13859__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09239_ _09241_/CLK line[39] VGND VGND VPWR VPWR _09240_/A sky130_fd_sc_hd__dfxtp_1
X_12250_ _12249_/Q _12257_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_11201_ _11191_/CLK line[40] VGND VGND VPWR VPWR _11202_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[4\].VALID\[4\].FF OVHB\[4\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[4\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10283__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _12177_/CLK line[104] VGND VGND VPWR VPWR _12182_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05377__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11132_ _11131_/Q _11137_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13594__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_MUX.MUX\[22\]_A2 _06543_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11063_ _11063_/CLK line[105] VGND VGND VPWR VPWR _11064_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08688__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07592__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10014_ _10013_/Q _10017_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06001__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DEC.DEC0.AND3_B A[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11965_ _11945_/CLK line[5] VGND VGND VPWR VPWR _11965_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11842__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13704_ _13703_/Q _13727_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_10916_ _10915_/Q _10927_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_11896_ _11895_/Q _11907_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05840__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13635_ _13631_/CLK line[15] VGND VGND VPWR VPWR _13635_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10458__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10847_ _10843_/CLK line[6] VGND VGND VPWR VPWR _10848_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[17\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13412__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13566_ _13565_/Q _13587_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_10778_ _10778_/A _10787_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13769__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12517_ _12523_/CLK line[1] VGND VGND VPWR VPWR _12517_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12673__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13131__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13497_ _13497_/CLK line[65] VGND VGND VPWR VPWR _13498_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07767__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12448_ _12447_/Q _12467_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06026__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10193__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12379_ _12387_/CLK line[66] VGND VGND VPWR VPWR _12379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[4\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _12430_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10921__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06940_ _06960_/CLK line[26] VGND VGND VPWR VPWR _06940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[2\].VALID\[6\].FF OVHB\[2\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[2\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06871_ _06870_/Q _06902_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13009__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08610_ _08610_/A _08617_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_05822_ _05836_/CLK line[27] VGND VGND VPWR VPWR _05822_/Q sky130_fd_sc_hd__dfxtp_1
X_09590_ _09590_/A _09597_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[5\].TOBUF OVHB\[12\].VALID\[5\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09072__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08541_ _08541_/CLK line[104] VGND VGND VPWR VPWR _08542_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13306__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05753_ _05753_/A _05782_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12848__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08472_ _08472_/A _08477_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_05684_ _05708_/CLK line[92] VGND VGND VPWR VPWR _05685_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05750__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07423_ _07393_/CLK line[105] VGND VGND VPWR VPWR _07423_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10368__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07354_ _07353_/Q _07357_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_06305_ _06305_/CLK _06306_/X VGND VGND VPWR VPWR _06285_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_109_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12583__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07285_ _07285_/CLK _07286_/X VGND VGND VPWR VPWR _07267_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07677__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09024_ _09023_/Q _09037_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06581__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06236_ _06272_/A wr VGND VGND VPWR VPWR _06236_/X sky130_fd_sc_hd__and2_1
XFILLER_102_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11199__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06167_ _06272_/A VGND VGND VPWR VPWR _06167_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10681__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09892__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05118_ _05122_/CLK line[80] VGND VGND VPWR VPWR _05118_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09247__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06098_ _06108_/CLK line[16] VGND VGND VPWR VPWR _06098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10831__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09926_ _09925_/Q _09947_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_05049_ _05048_/Q _05082_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[0\].FF OVHB\[30\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[30\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05925__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[12\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09857_ _09849_/CLK line[65] VGND VGND VPWR VPWR _09857_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[3\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _12045_/CLK sky130_fd_sc_hd__clkbuf_4
X_08808_ _08807_/Q _08827_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
X_09788_ _09787_/Q _09807_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04933__B1 A_h[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08739_ _08749_/CLK line[66] VGND VGND VPWR VPWR _08739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12758__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06756__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11750_ _11750_/A _11767_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[8\].FF OVHB\[0\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[0\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10707_/CLK line[67] VGND VGND VPWR VPWR _10702_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11691_/CLK line[3] VGND VGND VPWR VPWR _11681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10856__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13419_/Q _13447_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _10631_/Q _10647_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ _10571_/CLK line[4] VGND VGND VPWR VPWR _10564_/A sky130_fd_sc_hd__dfxtp_1
X_13351_ _13347_/CLK line[13] VGND VGND VPWR VPWR _13351_/Q sky130_fd_sc_hd__dfxtp_1
X_12302_ _12301_/Q _12327_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06491__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13282_ _13281_/Q _13307_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_10494_ _10493_/Q _10507_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12233_ _12227_/CLK line[14] VGND VGND VPWR VPWR _12233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12164_ _12164_/A _12187_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[23\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _09385_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[29\].VALID\[1\].FF OVHB\[29\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[29\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11115_ _11111_/CLK line[15] VGND VGND VPWR VPWR _11116_/A sky130_fd_sc_hd__dfxtp_1
X_12095_ _12109_/CLK line[79] VGND VGND VPWR VPWR _12095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09307__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11046_ _11046_/A _11067_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12997_ _12999_/CLK line[107] VGND VGND VPWR VPWR _12997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11572__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06666__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11948_ _11947_/Q _11977_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09042__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10188__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11879_ _11901_/CLK line[108] VGND VGND VPWR VPWR _11880_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08881__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13618_ _13598_/CLK line[121] VGND VGND VPWR VPWR _13618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13499__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[11\].TOBUF OVHB\[28\].VALID\[11\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_13549_ _13548_/Q _13552_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[1\].VALID\[14\].TOBUF OVHB\[1\].VALID\[14\].FF/Q OVHB\[1\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_07070_ _07069_/Q _07077_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13796__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06021_ _06023_/CLK line[104] VGND VGND VPWR VPWR _06022_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[15\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11747__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07972_ _07971_/Q _07987_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09217__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08121__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09711_ _09721_/CLK line[13] VGND VGND VPWR VPWR _09711_/Q sky130_fd_sc_hd__dfxtp_1
X_06923_ _06923_/CLK line[4] VGND VGND VPWR VPWR _06923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[22\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _09000_/CLK sky130_fd_sc_hd__clkbuf_4
X_09642_ _09641_/Q _09667_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06854_ _06853_/Q _06867_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12221__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[3\].FF OVHB\[27\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[27\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05805_ _05799_/CLK line[5] VGND VGND VPWR VPWR _05805_/Q sky130_fd_sc_hd__dfxtp_1
X_06785_ _06775_/CLK line[69] VGND VGND VPWR VPWR _06785_/Q sky130_fd_sc_hd__dfxtp_1
X_09573_ _09577_/CLK line[78] VGND VGND VPWR VPWR _09573_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[10\].TOBUF OVHB\[21\].VALID\[10\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05736_ _05736_/A _05747_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_08524_ _08524_/A _08547_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[4\]_A2 _13504_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05480__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[8\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ _08473_/CLK line[79] VGND VGND VPWR VPWR _08456_/A sky130_fd_sc_hd__dfxtp_1
X_05667_ _05671_/CLK line[70] VGND VGND VPWR VPWR _05668_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _07406_/A _07427_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08386_ _08385_/Q _08407_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[12\]_A1 _05020_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05598_ _05597_/Q _05607_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07337_ _07327_/CLK line[65] VGND VGND VPWR VPWR _07337_/Q sky130_fd_sc_hd__dfxtp_1
X_07268_ _07267_/Q _07287_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06219_ _06223_/CLK line[66] VGND VGND VPWR VPWR _06219_/Q sky130_fd_sc_hd__dfxtp_1
X_09007_ _09005_/CLK line[75] VGND VGND VPWR VPWR _09007_/Q sky130_fd_sc_hd__dfxtp_1
X_07199_ _07183_/CLK line[2] VGND VGND VPWR VPWR _07199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[6\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10561__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05655__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08031__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09909_ _09909_/A _09912_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13872__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12920_ _12920_/CLK _12921_/X VGND VGND VPWR VPWR _12902_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_74_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07870__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12488__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12851_ _12992_/A wr VGND VGND VPWR VPWR _12851_/X sky130_fd_sc_hd__and2_1
X_11802_ _11872_/A VGND VGND VPWR VPWR _11802_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[6\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[21\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _08615_/CLK sky130_fd_sc_hd__clkbuf_4
X_12782_ _12712_/A VGND VGND VPWR VPWR _12782_/Y sky130_fd_sc_hd__inv_2
XOVHB\[19\].VALID\[5\].TOBUF OVHB\[19\].VALID\[5\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _11757_/CLK line[32] VGND VGND VPWR VPWR _11733_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _05745_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09797__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[25\].VALID\[5\].FF OVHB\[25\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[25\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11664_ _11663_/Q _11697_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08056__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13402_/Q _13412_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _10627_/CLK line[42] VGND VGND VPWR VPWR _10615_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11595_ _11605_/CLK line[106] VGND VGND VPWR VPWR _11595_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13308_/CLK line[119] VGND VGND VPWR VPWR _13334_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08206__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10546_ _10545_/Q _10577_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12951__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13265_ _13265_/A _13272_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_10477_ _10473_/CLK line[107] VGND VGND VPWR VPWR _10477_/Q sky130_fd_sc_hd__dfxtp_1
X_12216_ _12204_/CLK line[120] VGND VGND VPWR VPWR _12216_/Q sky130_fd_sc_hd__dfxtp_1
X_13196_ _13194_/CLK line[56] VGND VGND VPWR VPWR _13197_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12147_ _12146_/Q _12152_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12078_ _12072_/CLK line[57] VGND VGND VPWR VPWR _12078_/Q sky130_fd_sc_hd__dfxtp_1
X_11029_ _11029_/A _11032_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07780__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12398__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06570_ _06570_/A _06587_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06396__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05521_ _05519_/CLK line[3] VGND VGND VPWR VPWR _05521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08240_ _08239_/Q _08267_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_05452_ _05451_/Q _05467_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08171_ _08175_/CLK line[77] VGND VGND VPWR VPWR _08172_/A sky130_fd_sc_hd__dfxtp_1
X_05383_ _05391_/CLK line[68] VGND VGND VPWR VPWR _05384_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[1\].TOBUF OVHB\[0\].VALID\[1\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07122_ _07121_/Q _07147_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[10\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _05360_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07020__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12861__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07053_ _07043_/CLK line[78] VGND VGND VPWR VPWR _07053_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[4\].TOBUF OVHB\[25\].VALID\[4\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07955__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[7\].FF OVHB\[23\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[23\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06004_ _06004_/A _06027_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11477__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07955_ _07981_/CLK line[106] VGND VGND VPWR VPWR _07956_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[13\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06906_ _06906_/A _06937_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08786__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07886_ _07885_/Q _07917_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09625_ _09625_/A _09632_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06837_ _06839_/CLK line[107] VGND VGND VPWR VPWR _06837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12886__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12101__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09556_ _09554_/CLK line[56] VGND VGND VPWR VPWR _09557_/A sky130_fd_sc_hd__dfxtp_1
X_06768_ _06767_/Q _06797_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08507_ _08507_/A _08512_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_05719_ _05739_/CLK line[108] VGND VGND VPWR VPWR _05719_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06699_ _06711_/CLK line[44] VGND VGND VPWR VPWR _06700_/A sky130_fd_sc_hd__dfxtp_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09487_ _09487_/A _09492_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _08410_/CLK line[57] VGND VGND VPWR VPWR _08438_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDECH.DEC0.AND0 A_h[7] A_h[8] VGND VGND VPWR VPWR _13990_/D sky130_fd_sc_hd__nor2_2
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[18\] _11435_/Z _13465_/Z _07095_/Z _13605_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[18] sky130_fd_sc_hd__mux4_1
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08369_ _08368_/Q _08372_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10400_ _10400_/CLK _10401_/X VGND VGND VPWR VPWR _10384_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11380_ _11380_/CLK _11381_/X VGND VGND VPWR VPWR _11370_/CLK sky130_fd_sc_hd__dlclkp_1
X_10331_ _13931_/X wr VGND VGND VPWR VPWR _10331_/X sky130_fd_sc_hd__and2_1
XFILLER_118_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10262_ _10192_/A VGND VGND VPWR VPWR _10262_/Y sky130_fd_sc_hd__inv_2
X_13050_ _13050_/CLK line[117] VGND VGND VPWR VPWR _13050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11387__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10291__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12001_ _12000_/Q _12012_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10193_ _10217_/CLK line[96] VGND VGND VPWR VPWR _10193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05385__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[31\].VALID\[3\].TOBUF OVHB\[31\].VALID\[3\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_13952_ _13950_/C _13950_/A _13950_/B _13957_/D VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__and4bb_4
XOVHB\[21\].VALID\[9\].FF OVHB\[21\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[21\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08696__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12903_ _12903_/A _12922_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_13883_ _13883_/A _13902_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12834_ _12820_/CLK line[18] VGND VGND VPWR VPWR _12835_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12764_/Q _12782_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11850__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11716_ _11706_/CLK line[19] VGND VGND VPWR VPWR _11716_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06944__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09320__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12708_/CLK line[83] VGND VGND VPWR VPWR _12696_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10466__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11647_ _11646_/Q _11662_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11578_ _11588_/CLK line[84] VGND VGND VPWR VPWR _11578_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13777__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13317_ _13316_/Q _13342_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_10529_ _10528_/Q _10542_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_13248_ _13254_/CLK line[94] VGND VGND VPWR VPWR _13248_/Q sky130_fd_sc_hd__dfxtp_1
X_13179_ _13178_/Q _13202_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05295__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07740_ _07740_/CLK _07741_/X VGND VGND VPWR VPWR _07724_/CLK sky130_fd_sc_hd__dlclkp_1
X_04952_ _04952_/A _04977_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07671_ _07672_/A wr VGND VGND VPWR VPWR _07671_/X sky130_fd_sc_hd__and2_1
XFILLER_19_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13017__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09410_ _09414_/CLK line[117] VGND VGND VPWR VPWR _09410_/Q sky130_fd_sc_hd__dfxtp_1
X_06622_ _06551_/A VGND VGND VPWR VPWR _06622_/Y sky130_fd_sc_hd__inv_2
XOVHB\[23\].VALID\[9\].TOBUF OVHB\[23\].VALID\[9\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09341_ _09340_/Q _09352_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_06553_ _06565_/CLK line[96] VGND VGND VPWR VPWR _06553_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05504_ _05503_/Q _05537_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_09272_ _09256_/CLK line[54] VGND VGND VPWR VPWR _09272_/Q sky130_fd_sc_hd__dfxtp_1
X_06484_ _06483_/Q _06517_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_05435_ _05445_/CLK line[106] VGND VGND VPWR VPWR _05436_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10376__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08223_ _08222_/Q _08232_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_08154_ _08134_/CLK line[55] VGND VGND VPWR VPWR _08154_/Q sky130_fd_sc_hd__dfxtp_1
X_05366_ _05365_/Q _05397_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_07105_ _07104_/Q _07112_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12591__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08085_ _08084_/Q _08092_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_05297_ _05299_/CLK line[43] VGND VGND VPWR VPWR _05297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07685__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07036_ _07030_/CLK line[56] VGND VGND VPWR VPWR _07036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08987_ _08986_/Q _09002_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07938_ _07946_/CLK line[84] VGND VGND VPWR VPWR _07938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05933__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07869_ _07868_/Q _07882_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09608_ _09626_/CLK line[94] VGND VGND VPWR VPWR _09608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10880_ _10872_/CLK line[21] VGND VGND VPWR VPWR _10880_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09539_ _09538_/Q _09562_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12766__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[4\].CGAND _13943_/X wr VGND VGND VPWR VPWR OVHB\[4\].CGAND/X sky130_fd_sc_hd__and2_4
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12560_/CLK line[31] VGND VGND VPWR VPWR _12550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _11500_/Q _11522_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12481_ _12480_/Q _12502_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _11440_/CLK line[17] VGND VGND VPWR VPWR _11432_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11363_ _11362_/Q _11382_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[1\].TOBUF OVHB\[7\].VALID\[1\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _13120_/CLK line[27] VGND VGND VPWR VPWR _13103_/A sky130_fd_sc_hd__dfxtp_1
X_10314_ _10314_/CLK line[18] VGND VGND VPWR VPWR _10314_/Q sky130_fd_sc_hd__dfxtp_1
X_11294_ _11302_/CLK line[82] VGND VGND VPWR VPWR _11294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[25\]_A0 _10329_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ _13032_/Q _13062_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12006__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10245_ _10245_/A _10262_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10176_ _10188_/CLK line[83] VGND VGND VPWR VPWR _10177_/A sky130_fd_sc_hd__dfxtp_1
X_13935_ _13933_/B _13934_/B _13934_/C _13934_/D VGND VGND VPWR VPWR _11872_/A sky130_fd_sc_hd__and4_4
XANTENNA_OVHB\[13\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13866_ _13907_/X wr VGND VGND VPWR VPWR _13866_/X sky130_fd_sc_hd__and2_1
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12817_ _12992_/A VGND VGND VPWR VPWR _12817_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13797_ _13907_/X VGND VGND VPWR VPWR _13797_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11580__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[16\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06674__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12748_ _12774_/CLK line[112] VGND VGND VPWR VPWR _12748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09050__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ _12678_/Q _12712_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09985__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06971__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05220_ _05220_/CLK _05221_/X VGND VGND VPWR VPWR _05214_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[23\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[14\].TOBUF OVHB\[14\].VALID\[14\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_05151_ _05152_/A wr VGND VGND VPWR VPWR _05151_/X sky130_fd_sc_hd__and2_1
X_05082_ _05152_/A VGND VGND VPWR VPWR _05082_/Y sky130_fd_sc_hd__inv_2
X_08910_ _08922_/CLK line[31] VGND VGND VPWR VPWR _08910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09890_ _09908_/CLK line[95] VGND VGND VPWR VPWR _09890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08841_ _08841_/A _08862_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11755__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06849__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08772_ _08762_/CLK line[81] VGND VGND VPWR VPWR _08772_/Q sky130_fd_sc_hd__dfxtp_1
X_05984_ _05984_/CLK line[87] VGND VGND VPWR VPWR _05984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09225__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07723_ _07723_/A _07742_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_04935_ A_h[17] _04935_/B2 A_h[17] _04935_/B2 VGND VGND VPWR VPWR _04935_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07654_ _07644_/CLK line[82] VGND VGND VPWR VPWR _07654_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06605_ _06604_/Q _06622_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11490__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07585_ _07584_/Q _07602_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09324_ _09320_/CLK line[92] VGND VGND VPWR VPWR _09324_/Q sky130_fd_sc_hd__dfxtp_1
X_06536_ _06528_/CLK line[83] VGND VGND VPWR VPWR _06536_/Q sky130_fd_sc_hd__dfxtp_1
X_09255_ _09254_/Q _09282_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_06467_ _06466_/Q _06482_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _08300_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08206_ _08208_/CLK line[93] VGND VGND VPWR VPWR _08206_/Q sky130_fd_sc_hd__dfxtp_1
X_05418_ _05424_/CLK line[84] VGND VGND VPWR VPWR _05418_/Q sky130_fd_sc_hd__dfxtp_1
X_06398_ _06408_/CLK line[20] VGND VGND VPWR VPWR _06399_/A sky130_fd_sc_hd__dfxtp_1
X_09186_ _09200_/CLK line[29] VGND VGND VPWR VPWR _09187_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05349_ _05349_/A _05362_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_08137_ _08136_/Q _08162_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[15\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08068_ _08070_/CLK line[30] VGND VGND VPWR VPWR _08068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07019_ _07018_/Q _07042_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10030_ _10042_/CLK line[31] VGND VGND VPWR VPWR _10030_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11665__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05663__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[31\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _11870_/CLK sky130_fd_sc_hd__clkbuf_4
X_11981_ _11981_/A _12012_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13880__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[25\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[4\].CGAND_A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13720_ _13719_/Q _13727_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08974__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10932_ _10930_/CLK line[59] VGND VGND VPWR VPWR _10932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[5\].VALID\[6\].TOBUF OVHB\[5\].VALID\[6\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_13651_ _13631_/CLK line[8] VGND VGND VPWR VPWR _13651_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12496__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10863_ _10862_/Q _10892_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_12602_ _12602_/A _12607_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _13581_/Q _13587_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_10794_ _10804_/CLK line[124] VGND VGND VPWR VPWR _10794_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12533_ _12523_/CLK line[9] VGND VGND VPWR VPWR _12534_/A sky130_fd_sc_hd__dfxtp_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ _12463_/Q _12467_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _11415_/CLK _11416_/X VGND VGND VPWR VPWR _11395_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10744__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12395_ _12395_/CLK _12396_/X VGND VGND VPWR VPWR _12387_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13120__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05838__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _05115_/CLK sky130_fd_sc_hd__clkbuf_4
X_11346_ _11311_/A wr VGND VGND VPWR VPWR _11346_/X sky130_fd_sc_hd__and2_1
XANTENNA__08214__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11277_ _11311_/A VGND VGND VPWR VPWR _11277_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08511__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13016_ _13015_/Q _13027_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_10228_ _10248_/CLK line[112] VGND VGND VPWR VPWR _10228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10159_ _10158_/Q _10192_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05573__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ _13923_/C _13923_/B _13922_/B _13923_/D VGND VGND VPWR VPWR _13918_/X sky130_fd_sc_hd__and4bb_4
XFILLER_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13849_ _13845_/CLK line[98] VGND VGND VPWR VPWR _13849_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10919__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _11485_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07370_ _07380_/CLK line[95] VGND VGND VPWR VPWR _07370_/Q sky130_fd_sc_hd__dfxtp_1
X_06321_ _06320_/Q _06342_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_09040_ _09068_/CLK line[90] VGND VGND VPWR VPWR _09041_/A sky130_fd_sc_hd__dfxtp_1
X_06252_ _06244_/CLK line[81] VGND VGND VPWR VPWR _06252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05203_ _05202_/Q _05222_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10654__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06183_ _06182_/Q _06202_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[9\].VALID\[7\].FF OVHB\[9\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[9\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[1\].TOBUF OVHB\[12\].VALID\[1\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13030__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05748__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05134_ _05122_/CLK line[82] VGND VGND VPWR VPWR _05135_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09942_ _09942_/A _09947_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_05065_ _05064_/Q _05082_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07963__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09873_ _09849_/CLK line[73] VGND VGND VPWR VPWR _09873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08824_ _08824_/A _08827_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06579__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08755_ _08755_/CLK _08756_/X VGND VGND VPWR VPWR _08749_/CLK sky130_fd_sc_hd__dlclkp_1
X_05967_ _05966_/Q _05992_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[7\]_A0 _11410_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07706_ _07672_/A wr VGND VGND VPWR VPWR _07706_/X sky130_fd_sc_hd__and2_1
X_04918_ _04917_/Y _04918_/A2 _04915_/Y _04918_/B2 VGND VGND VPWR VPWR _04918_/Y sky130_fd_sc_hd__a22oi_4
X_08686_ _13922_/X wr VGND VGND VPWR VPWR _08686_/X sky130_fd_sc_hd__and2_1
X_05898_ _05902_/CLK line[62] VGND VGND VPWR VPWR _05898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07637_ _07672_/A VGND VGND VPWR VPWR _07637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10829__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13205__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07568_ _07572_/CLK line[48] VGND VGND VPWR VPWR _07568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07203__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09307_ _09307_/CLK line[70] VGND VGND VPWR VPWR _09307_/Q sky130_fd_sc_hd__dfxtp_1
X_06519_ _06518_/Q _06552_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_07499_ _07498_/Q _07532_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_09238_ _09237_/Q _09247_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_09169_ _09147_/CLK line[7] VGND VGND VPWR VPWR _09169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11200_ _11200_/A _11207_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_12180_ _12180_/A _12187_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11131_ _11111_/CLK line[8] VGND VGND VPWR VPWR _11131_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[30\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11062_ _11062_/A _11067_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[22\]_A3 _13613_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06132__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[7\].VALID\[9\].FF OVHB\[7\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[7\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11395__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10013_ _10011_/CLK line[9] VGND VGND VPWR VPWR _10013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06489__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05393__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _11964_/A _11977_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_13703_ _13701_/CLK line[46] VGND VGND VPWR VPWR _13703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10915_ _10903_/CLK line[37] VGND VGND VPWR VPWR _10915_/Q sky130_fd_sc_hd__dfxtp_1
X_11895_ _11901_/CLK line[101] VGND VGND VPWR VPWR _11895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[11\].TOBUF OVHB\[8\].VALID\[11\].FF/Q OVHB\[8\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_13634_ _13633_/Q _13657_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_10846_ _10845_/Q _10857_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07113__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[23\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13565_ _13559_/CLK line[111] VGND VGND VPWR VPWR _13565_/Q sky130_fd_sc_hd__dfxtp_1
X_10777_ _10783_/CLK line[102] VGND VGND VPWR VPWR _10778_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12516_ _12515_/Q _12537_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06952__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06307__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13496_ _13495_/Q _13517_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_12447_ _12449_/CLK line[97] VGND VGND VPWR VPWR _12447_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06026__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05568__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ _12377_/Q _12397_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13785__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11329_ _11343_/CLK line[98] VGND VGND VPWR VPWR _11330_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08879__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06870_ _06892_/CLK line[122] VGND VGND VPWR VPWR _06870_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[10\].TOBUF OVHB\[1\].VALID\[10\].FF/Q OVHB\[1\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_05821_ _05820_/Q _05852_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08540_ _08539_/Q _08547_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_05752_ _05756_/CLK line[123] VGND VGND VPWR VPWR _05753_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[10\].VALID\[6\].TOBUF OVHB\[10\].VALID\[6\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__09503__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08471_ _08473_/CLK line[72] VGND VGND VPWR VPWR _08472_/A sky130_fd_sc_hd__dfxtp_1
X_05683_ _05682_/Q _05712_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_07422_ _07421_/Q _07427_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08119__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[8\].V OVHB\[8\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[8\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07601__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07353_ _07327_/CLK line[73] VGND VGND VPWR VPWR _07353_/Q sky130_fd_sc_hd__dfxtp_1
X_06304_ _06303_/Q _06307_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_07284_ _07283_/Q _07287_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10384__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09023_ _09005_/CLK line[68] VGND VGND VPWR VPWR _09023_/Q sky130_fd_sc_hd__dfxtp_1
X_06235_ _06235_/CLK _06236_/X VGND VGND VPWR VPWR _06223_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10962__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05478__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06166_ _06272_/A wr VGND VGND VPWR VPWR _06166_/X sky130_fd_sc_hd__and2_1
XANTENNA__10681__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13695__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[23\].VALID\[14\].FF OVHB\[23\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[23\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05117_ _05152_/A VGND VGND VPWR VPWR _05117_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06097_ _06272_/A VGND VGND VPWR VPWR _06097_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07693__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09925_ _09925_/CLK line[111] VGND VGND VPWR VPWR _09925_/Q sky130_fd_sc_hd__dfxtp_1
X_05048_ _05058_/CLK line[48] VGND VGND VPWR VPWR _05048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09856_ _09855_/Q _09877_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].V OVHB\[31\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[31\].V/Q sky130_fd_sc_hd__dfrtp_1
XOVHB\[16\].VALID\[1\].FF OVHB\[16\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[16\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08807_ _08823_/CLK line[97] VGND VGND VPWR VPWR _08807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06102__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09787_ _09793_/CLK line[33] VGND VGND VPWR VPWR _09787_/Q sky130_fd_sc_hd__dfxtp_1
X_06999_ _07001_/CLK line[39] VGND VGND VPWR VPWR _06999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11943__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08738_ _08738_/A _08757_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04933__B2 _04933_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05941__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10559__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ _08663_/CLK line[34] VGND VGND VPWR VPWR _08670_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10699_/Q _10717_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11679_/Q _11697_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _10627_/CLK line[35] VGND VGND VPWR VPWR _10631_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12774__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13350_ _13349_/Q _13377_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_10562_ _10561_/Q _10577_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12301_ _12311_/CLK line[45] VGND VGND VPWR VPWR _12301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13281_ _13285_/CLK line[109] VGND VGND VPWR VPWR _13281_/Q sky130_fd_sc_hd__dfxtp_1
X_10493_ _10473_/CLK line[100] VGND VGND VPWR VPWR _10493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _12232_/A _12257_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[31\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12163_ _12177_/CLK line[110] VGND VGND VPWR VPWR _12164_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[1\].TOBUF OVHB\[19\].VALID\[1\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_11114_ _11113_/Q _11137_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_12094_ _12093_/Q _12117_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11045_ _11063_/CLK line[111] VGND VGND VPWR VPWR _11046_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06797__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].V OVHB\[22\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[22\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07108__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12949__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ _12995_/Q _13027_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[24\].VALID\[12\].TOBUF OVHB\[24\].VALID\[12\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_11947_ _11945_/CLK line[11] VGND VGND VPWR VPWR _11947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[3\].FF OVHB\[14\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[14\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11878_ _11878_/A _11907_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_13617_ _13616_/Q _13622_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12684__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10829_ _10843_/CLK line[12] VGND VGND VPWR VPWR _10829_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[7\].FF OVHB\[31\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[31\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07778__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06682__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13548_ _13528_/CLK line[89] VGND VGND VPWR VPWR _13548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[7\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13479_ _13478_/Q _13482_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09993__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06020_ _06020_/A _06027_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[21\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10932__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07971_ _07981_/CLK line[99] VGND VGND VPWR VPWR _07971_/Q sky130_fd_sc_hd__dfxtp_1
X_09710_ _09709_/Q _09737_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_06922_ _06922_/A _06937_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12502__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07018__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].V OVHB\[13\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[13\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09641_ _09659_/CLK line[109] VGND VGND VPWR VPWR _09641_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12859__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06853_ _06839_/CLK line[100] VGND VGND VPWR VPWR _06853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11763__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12221__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05804_ _05803_/Q _05817_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06857__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09572_ _09572_/A _09597_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
X_06784_ _06783_/Q _06797_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[0\].TOBUF OVHB\[25\].VALID\[0\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09233__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08523_ _08541_/CLK line[110] VGND VGND VPWR VPWR _08524_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05116__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05735_ _05739_/CLK line[101] VGND VGND VPWR VPWR _05736_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[4\]_A3 _06854_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ _08454_/A _08477_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05666_ _05666_/A _05677_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_07405_ _07393_/CLK line[111] VGND VGND VPWR VPWR _07406_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08385_ _08383_/CLK line[47] VGND VGND VPWR VPWR _08385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[12\]_A2 _13490_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05597_ _05575_/CLK line[38] VGND VGND VPWR VPWR _05597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06592__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07336_ _07335_/Q _07357_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07267_ _07267_/CLK line[33] VGND VGND VPWR VPWR _07267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09006_ _09005_/Q _09037_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[5\].FF OVHB\[12\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[12\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06218_ _06218_/A _06237_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08162__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07198_ _07197_/Q _07217_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11938__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06149_ _06147_/CLK line[34] VGND VGND VPWR VPWR _06149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09408__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09908_ _09908_/CLK line[89] VGND VGND VPWR VPWR _09909_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09839_ _09839_/A _09842_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11673__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06767__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _12850_/CLK _12851_/X VGND VGND VPWR VPWR _12820_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_100_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05671__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09143__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11801_ _11872_/A wr VGND VGND VPWR VPWR _11801_/X sky130_fd_sc_hd__and2_1
XFILLER_15_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10289__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12781_ _12712_/A wr VGND VGND VPWR VPWR _12781_/X sky130_fd_sc_hd__and2_1
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08982__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11732_ _11872_/A VGND VGND VPWR VPWR _11732_/Y sky130_fd_sc_hd__inv_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08337__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[6\].TOBUF OVHB\[17\].VALID\[6\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11691_/CLK line[0] VGND VGND VPWR VPWR _11663_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07598__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08056__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ _13394_/CLK line[22] VGND VGND VPWR VPWR _13402_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ _10613_/Q _10647_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _11593_/Q _11627_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13333_ _13332_/Q _13342_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10545_ _10571_/CLK line[10] VGND VGND VPWR VPWR _10545_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06007__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13264_ _13254_/CLK line[87] VGND VGND VPWR VPWR _13265_/A sky130_fd_sc_hd__dfxtp_1
X_10476_ _10475_/Q _10507_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11848__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12215_ _12214_/Q _12222_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13195_ _13195_/A _13202_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05846__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09318__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08222__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12146_ _12130_/CLK line[88] VGND VGND VPWR VPWR _12146_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04939__A2_N _04939_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ _12076_/Q _12082_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[7\].FF OVHB\[10\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[10\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11028_ _11002_/CLK line[89] VGND VGND VPWR VPWR _11029_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05581__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09631__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10199__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12979_ _12978_/Q _12992_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
X_05520_ _05519_/Q _05537_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05451_ _05445_/CLK line[99] VGND VGND VPWR VPWR _05451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12992__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13303__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _08169_/Q _08197_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_05382_ _05381_/Q _05397_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_07121_ _07117_/CLK line[109] VGND VGND VPWR VPWR _07121_/Q sky130_fd_sc_hd__dfxtp_1
X_07052_ _07051_/Q _07077_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[5\].TOBUF OVHB\[23\].VALID\[5\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_127_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06003_ _06023_/CLK line[110] VGND VGND VPWR VPWR _06004_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10662__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10017__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05756__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09806__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08132__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07954_ _07953_/Q _07987_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07971__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06905_ _06923_/CLK line[10] VGND VGND VPWR VPWR _06906_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12589__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07885_ _07905_/CLK line[74] VGND VGND VPWR VPWR _07885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09624_ _09626_/CLK line[87] VGND VGND VPWR VPWR _09625_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06836_ _06835_/Q _06867_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12886__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09555_ _09554_/Q _09562_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_06767_ _06775_/CLK line[75] VGND VGND VPWR VPWR _06767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09898__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08506_ _08480_/CLK line[88] VGND VGND VPWR VPWR _08507_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05718_ _05717_/Q _05747_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ _09482_/CLK line[24] VGND VGND VPWR VPWR _09487_/A sky130_fd_sc_hd__dfxtp_1
X_06698_ _06697_/Q _06727_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08437_ _08436_/Q _08442_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10837__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05649_ _05671_/CLK line[76] VGND VGND VPWR VPWR _05650_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDECH.DEC0.AND1 A_h[8] A_h[7] VGND VGND VPWR VPWR _13957_/D sky130_fd_sc_hd__and2b_2
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08307__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08368_ _08358_/CLK line[25] VGND VGND VPWR VPWR _08368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07211__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07319_ _07318_/Q _07322_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_08299_ _08298_/Q _08302_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11311__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10330_ _10330_/CLK _10331_/X VGND VGND VPWR VPWR _10314_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_3_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ _10192_/A wr VGND VGND VPWR VPWR _10261_/X sky130_fd_sc_hd__and2_1
XANTENNA__09138__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ _12002_/CLK line[21] VGND VGND VPWR VPWR _12000_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].CGAND _05152_/A wr VGND VGND VPWR VPWR OVHB\[0\].CG/GATE sky130_fd_sc_hd__and2_4
X_10192_ _10192_/A VGND VGND VPWR VPWR _10192_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13951_ _13950_/C _13950_/B _13950_/A _13957_/D VGND VGND VPWR VPWR _13951_/X sky130_fd_sc_hd__and4bb_4
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12902_ _12902_/CLK line[49] VGND VGND VPWR VPWR _12903_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06497__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13882_ _13882_/CLK line[113] VGND VGND VPWR VPWR _13883_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12833_ _12832_/Q _12852_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12764_ _12774_/CLK line[114] VGND VGND VPWR VPWR _12764_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11715_ _11715_/A _11732_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12695_ _12694_/Q _12712_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[3\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11646_ _11636_/CLK line[115] VGND VGND VPWR VPWR _11646_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07121__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12962__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _11576_/Q _11592_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13308_/CLK line[125] VGND VGND VPWR VPWR _13316_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06960__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10528_ _10520_/CLK line[116] VGND VGND VPWR VPWR _10528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11578__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13247_ _13246_/Q _13272_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_10459_ _10459_/A _10472_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09048__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ _13194_/CLK line[62] VGND VGND VPWR VPWR _13178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13793__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12128_/Q _12152_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08887__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07146__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04951_ _04947_/CLK line[13] VGND VGND VPWR VPWR _04952_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[0\].FF OVHB\[3\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[3\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[14\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12202__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07670_ _07670_/CLK _07671_/X VGND VGND VPWR VPWR _07644_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[14\].VALID\[10\].TOBUF OVHB\[14\].VALID\[10\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_38_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06621_ _06551_/A wr VGND VGND VPWR VPWR _06621_/X sky130_fd_sc_hd__and2_1
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09340_ _09320_/CLK line[85] VGND VGND VPWR VPWR _09340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06552_ _06551_/A VGND VGND VPWR VPWR _06552_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09511__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05503_ _05519_/CLK line[0] VGND VGND VPWR VPWR _05503_/Q sky130_fd_sc_hd__dfxtp_1
X_09271_ _09270_/Q _09282_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_06483_ _06489_/CLK line[64] VGND VGND VPWR VPWR _06483_/Q sky130_fd_sc_hd__dfxtp_1
X_08222_ _08208_/CLK line[86] VGND VGND VPWR VPWR _08222_/Q sky130_fd_sc_hd__dfxtp_1
X_05434_ _05433_/Q _05467_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[14\].FF OVHB\[28\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[28\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08153_ _08152_/Q _08162_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_05365_ _05391_/CLK line[74] VGND VGND VPWR VPWR _05365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07104_ _07098_/CLK line[87] VGND VGND VPWR VPWR _07104_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06870__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[7\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08084_ _08070_/CLK line[23] VGND VGND VPWR VPWR _08084_/Q sky130_fd_sc_hd__dfxtp_1
X_05296_ _05295_/Q _05327_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11488__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10392__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07035_ _07035_/A _07042_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05486__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08797__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08986_ _08972_/CLK line[51] VGND VGND VPWR VPWR _08986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07937_ _07937_/A _07952_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07868_ _07854_/CLK line[52] VGND VGND VPWR VPWR _07868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06110__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09607_ _09606_/Q _09632_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06819_ _06818_/Q _06832_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11951__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07799_ _07798_/Q _07812_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_09538_ _09554_/CLK line[62] VGND VGND VPWR VPWR _09538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[30\] _09469_/Z _13459_/Z _09609_/Z _13599_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[30] sky130_fd_sc_hd__mux4_1
XOVHB\[1\].VALID\[2\].FF OVHB\[1\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[1\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10567__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09469_ _09468_/Q _09492_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _11500_/CLK line[63] VGND VGND VPWR VPWR _11500_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12490_/CLK line[127] VGND VGND VPWR VPWR _12480_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08037__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13878__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _11430_/Q _11452_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07876__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11362_ _11370_/CLK line[113] VGND VGND VPWR VPWR _11362_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13101_ _13100_/Q _13132_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11976__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10313_ _10312_/Q _10332_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_11293_ _11292_/Q _11312_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[2\].TOBUF OVHB\[5\].VALID\[2\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[25\]_A1 _07039_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13032_ _13050_/CLK line[123] VGND VGND VPWR VPWR _13032_/Q sky130_fd_sc_hd__dfxtp_1
X_10244_ _10248_/CLK line[114] VGND VGND VPWR VPWR _10245_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10175_ _10174_/Q _10192_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08500__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13118__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13934_ _13933_/B _13934_/B _13934_/C _13934_/D VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__and4b_4
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[5\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13865_ _13865_/CLK _13866_/X VGND VGND VPWR VPWR _13845_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12816_ _12992_/A wr VGND VGND VPWR VPWR _12816_/X sky130_fd_sc_hd__and2_1
XFILLER_43_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13796_ _13907_/X wr VGND VGND VPWR VPWR _13796_/X sky130_fd_sc_hd__and2_1
XFILLER_62_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10477__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12747_ _12712_/A VGND VGND VPWR VPWR _12747_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12708_/CLK line[80] VGND VGND VPWR VPWR _12678_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11629_ _11628_/Q _11662_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12692__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12047__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07786__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05150_ _05150_/CLK _05151_/X VGND VGND VPWR VPWR _05122_/CLK sky130_fd_sc_hd__dlclkp_1
X_05081_ _05152_/A wr VGND VGND VPWR VPWR _05081_/X sky130_fd_sc_hd__and2_1
XFILLER_98_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10940__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08840_ _08850_/CLK line[127] VGND VGND VPWR VPWR _08841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08410__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[14\].FF OVHB\[0\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[0\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08771_ _08770_/Q _08792_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05983_ _05982_/Q _05992_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13028__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07722_ _07724_/CLK line[113] VGND VGND VPWR VPWR _07723_/A sky130_fd_sc_hd__dfxtp_1
X_04934_ A_h[19] _04934_/B2 A_h[19] _04934_/B2 VGND VGND VPWR VPWR _04936_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07026__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12867__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07653_ _07653_/A _07672_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06604_ _06596_/CLK line[114] VGND VGND VPWR VPWR _06604_/Q sky130_fd_sc_hd__dfxtp_1
X_07584_ _07572_/CLK line[50] VGND VGND VPWR VPWR _07584_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09241__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09323_ _09322_/Q _09352_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_06535_ _06534_/Q _06552_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[12\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13341__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09254_ _09256_/CLK line[60] VGND VGND VPWR VPWR _09254_/Q sky130_fd_sc_hd__dfxtp_1
X_06466_ _06464_/CLK line[51] VGND VGND VPWR VPWR _06466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08205_ _08204_/Q _08232_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_05417_ _05416_/Q _05432_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_09185_ _09184_/Q _09212_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_06397_ _06396_/Q _06412_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08136_ _08134_/CLK line[61] VGND VGND VPWR VPWR _08136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05348_ _05332_/CLK line[52] VGND VGND VPWR VPWR _05349_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12107__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08067_ _08066_/Q _08092_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05279_ _05278_/Q _05292_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07018_ _07030_/CLK line[62] VGND VGND VPWR VPWR _07018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[5\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09416__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08969_ _08969_/A _09002_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13516__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ _12002_/CLK line[26] VGND VGND VPWR VPWR _11981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10931_ _10930_/Q _10962_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[31\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[4\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[12\].FF OVHB\[24\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[24\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[23\].CGAND_A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11681__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06775__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _13650_/A _13657_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10862_ _10872_/CLK line[27] VGND VGND VPWR VPWR _10862_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09151__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[7\].TOBUF OVHB\[3\].VALID\[7\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[8\].CGAND_A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12601_ _12601_/CLK line[40] VGND VGND VPWR VPWR _12602_/A sky130_fd_sc_hd__dfxtp_1
X_13581_ _13559_/CLK line[104] VGND VGND VPWR VPWR _13581_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _10792_/Q _10822_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08990__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12532_ _12531_/Q _12537_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12463_ _12449_/CLK line[105] VGND VGND VPWR VPWR _12463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11414_ _11413_/Q _11417_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_12394_ _12393_/Q _12397_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_11345_ _11345_/CLK _11346_/X VGND VGND VPWR VPWR _11343_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12017__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06015__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09176__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11276_ _11311_/A wr VGND VGND VPWR VPWR _11276_/X sky130_fd_sc_hd__and2_1
XANTENNA__11856__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[14\].FF OVHB\[14\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[14\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13015_ _12999_/CLK line[101] VGND VGND VPWR VPWR _13015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10227_ _10192_/A VGND VGND VPWR VPWR _10227_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09326__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _10188_/CLK line[80] VGND VGND VPWR VPWR _10158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10089_ _10088_/Q _10122_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_13917_ _13922_/B _13923_/B _13923_/C _13923_/D VGND VGND VPWR VPWR _07111_/A sky130_fd_sc_hd__nor4b_4
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _13847_/Q _13867_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13779_ _13763_/CLK line[66] VGND VGND VPWR VPWR _13779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06320_ _06320_/CLK line[127] VGND VGND VPWR VPWR _06320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06251_ _06250_/Q _06272_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _10855_/CLK sky130_fd_sc_hd__clkbuf_4
X_05202_ _05214_/CLK line[113] VGND VGND VPWR VPWR _05202_/Q sky130_fd_sc_hd__dfxtp_1
X_06182_ _06186_/CLK line[49] VGND VGND VPWR VPWR _06182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[10\].VALID\[2\].TOBUF OVHB\[10\].VALID\[2\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[19\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _07985_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[14\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05133_ _05132_/Q _05152_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[1\].FF OVHB\[24\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[24\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09941_ _09925_/CLK line[104] VGND VGND VPWR VPWR _09942_/A sky130_fd_sc_hd__dfxtp_1
X_05064_ _05058_/CLK line[50] VGND VGND VPWR VPWR _05064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10670__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09872_ _09871_/Q _09877_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05764__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08140__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08823_ _08823_/CLK line[105] VGND VGND VPWR VPWR _08824_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08754_ _08754_/A _08757_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_05966_ _05984_/CLK line[93] VGND VGND VPWR VPWR _05966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07705_ _07705_/CLK _07706_/X VGND VGND VPWR VPWR _07679_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.MUX\[7\]_A1 _05600_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04917_ A_h[16] VGND VGND VPWR VPWR _04917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12597__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08685_ _08685_/CLK _08686_/X VGND VGND VPWR VPWR _08663_/CLK sky130_fd_sc_hd__dlclkp_1
X_05897_ _05896_/Q _05922_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07636_ _07672_/A wr VGND VGND VPWR VPWR _07636_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.MUX\[15\]_A0 _11396_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07567_ _07672_/A VGND VGND VPWR VPWR _07567_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11006__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09306_ _09305_/Q _09317_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06518_ _06528_/CLK line[80] VGND VGND VPWR VPWR _06518_/Q sky130_fd_sc_hd__dfxtp_1
X_07498_ _07518_/CLK line[16] VGND VGND VPWR VPWR _07498_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05004__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09237_ _09241_/CLK line[38] VGND VGND VPWR VPWR _09237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10845__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06449_ _06449_/A _06482_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13221__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05939__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08315__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09168_ _09168_/A _09177_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[10\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08119_ _08113_/CLK line[39] VGND VGND VPWR VPWR _08119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09099_ _09085_/CLK line[103] VGND VGND VPWR VPWR _09099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11130_ _11130_/A _11137_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[30\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10580__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11061_ _11063_/CLK line[104] VGND VGND VPWR VPWR _11062_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[18\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _07600_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[15\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10012_ _10011_/Q _10017_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[4\].VALID\[12\].TOBUF OVHB\[4\].VALID\[12\].FF/Q OVHB\[4\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_64_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[3\].FF OVHB\[22\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[22\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11963_ _11945_/CLK line[4] VGND VGND VPWR VPWR _11964_/A sky130_fd_sc_hd__dfxtp_1
X_13702_ _13702_/A _13727_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[3\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10914_ _10913_/Q _10927_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_11894_ _11894_/A _11907_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_13633_ _13631_/CLK line[14] VGND VGND VPWR VPWR _13633_/Q sky130_fd_sc_hd__dfxtp_1
X_10845_ _10843_/CLK line[5] VGND VGND VPWR VPWR _10845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10776_ _10775_/Q _10787_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_13564_ _13564_/A _13587_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10755__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12515_ _12523_/CLK line[15] VGND VGND VPWR VPWR _12515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13495_ _13497_/CLK line[79] VGND VGND VPWR VPWR _13495_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[27\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12446_ _12445_/Q _12467_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12970__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12377_ _12387_/CLK line[65] VGND VGND VPWR VPWR _12377_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11328_ _11327_/Q _11347_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11586__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11259_ _11251_/CLK line[66] VGND VGND VPWR VPWR _11260_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[10\].FF OVHB\[20\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[20\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09056__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05820_ _05836_/CLK line[26] VGND VGND VPWR VPWR _05820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _07215_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_48_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05751_ _05750_/Q _05782_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12210__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08470_ _08469_/Q _08477_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_05682_ _05708_/CLK line[91] VGND VGND VPWR VPWR _05682_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07304__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07421_ _07393_/CLK line[104] VGND VGND VPWR VPWR _07421_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[5\].FF OVHB\[20\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[20\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07601__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07352_ _07351_/Q _07357_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_06303_ _06285_/CLK line[105] VGND VGND VPWR VPWR _06303_/Q sky130_fd_sc_hd__dfxtp_1
X_07283_ _07267_/CLK line[41] VGND VGND VPWR VPWR _07283_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[12\].FF OVHB\[10\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[10\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09022_ _09022_/A _09037_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_06234_ _06233_/Q _06237_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06165_ _06165_/CLK _06166_/X VGND VGND VPWR VPWR _06147_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_85_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05116_ _05152_/A wr VGND VGND VPWR VPWR _05116_/X sky130_fd_sc_hd__and2_1
X_06096_ _06272_/A wr VGND VGND VPWR VPWR _06096_/X sky130_fd_sc_hd__and2_1
XANTENNA__11496__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09924_ _09924_/A _09947_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_05047_ _05152_/A VGND VGND VPWR VPWR _05047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05494__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09855_ _09849_/CLK line[79] VGND VGND VPWR VPWR _09855_/Q sky130_fd_sc_hd__dfxtp_1
X_08806_ _08805_/Q _08827_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09786_ _09785_/Q _09807_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_06998_ _06997_/Q _07007_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05949_ _05929_/CLK line[71] VGND VGND VPWR VPWR _05950_/A sky130_fd_sc_hd__dfxtp_1
X_08737_ _08749_/CLK line[65] VGND VGND VPWR VPWR _08738_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12120__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[14\].TOBUF OVHB\[27\].VALID\[14\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_08668_ _08667_/Q _08687_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[6\].FF OVHB\[19\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[19\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _07633_/CLK line[66] VGND VGND VPWR VPWR _07619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08599_ _08609_/CLK line[2] VGND VGND VPWR VPWR _08600_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[28\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10629_/Q _10647_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _10571_/CLK line[3] VGND VGND VPWR VPWR _10561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _12299_/Q _12327_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05669__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13280_ _13279_/Q _13307_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08045__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10492_ _10491_/Q _10507_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13886__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12231_ _12227_/CLK line[13] VGND VGND VPWR VPWR _12232_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12162_ _12161_/Q _12187_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11113_ _11111_/CLK line[14] VGND VGND VPWR VPWR _11113_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[2\].TOBUF OVHB\[17\].VALID\[2\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12093_ _12109_/CLK line[78] VGND VGND VPWR VPWR _12093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11044_ _11043_/Q _11067_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[13\].TOBUF OVHB\[20\].VALID\[13\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09604__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12995_ _12999_/CLK line[106] VGND VGND VPWR VPWR _12995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13126__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11946_ _11946_/A _11977_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11877_ _11901_/CLK line[107] VGND VGND VPWR VPWR _11878_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XMUX.MUX\[5\] _10846_/Z _05036_/Z _13506_/Z _05176_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[5] sky130_fd_sc_hd__mux4_1
X_13616_ _13598_/CLK line[120] VGND VGND VPWR VPWR _13616_/Q sky130_fd_sc_hd__dfxtp_1
X_10828_ _10827_/Q _10857_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05222__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10485__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13547_ _13546_/Q _13552_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
X_10759_ _10783_/CLK line[108] VGND VGND VPWR VPWR _10759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05579__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13478_ _13468_/CLK line[57] VGND VGND VPWR VPWR _13478_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[8\].FF OVHB\[17\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[17\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12429_ _12428_/Q _12432_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07794__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[14\].FF OVHB\[5\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[5\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07970_ _07970_/A _07987_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06203__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06921_ _06923_/CLK line[3] VGND VGND VPWR VPWR _06922_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].INV _13964_/X VGND VGND VPWR VPWR OVHB\[19\].INV/Y sky130_fd_sc_hd__inv_2
X_09640_ _09639_/Q _09667_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_06852_ _06851_/Q _06867_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05803_ _05799_/CLK line[4] VGND VGND VPWR VPWR _05803_/Q sky130_fd_sc_hd__dfxtp_1
X_09571_ _09577_/CLK line[77] VGND VGND VPWR VPWR _09572_/A sky130_fd_sc_hd__dfxtp_1
X_06783_ _06775_/CLK line[68] VGND VGND VPWR VPWR _06783_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13036__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08522_ _08521_/Q _08547_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_05734_ _05734_/A _05747_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05116__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[1\].TOBUF OVHB\[23\].VALID\[1\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07034__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12875__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08453_ _08473_/CLK line[78] VGND VGND VPWR VPWR _08454_/A sky130_fd_sc_hd__dfxtp_1
X_05665_ _05671_/CLK line[69] VGND VGND VPWR VPWR _05666_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07404_ _07404_/A _07427_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07969__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[20\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08384_ _08384_/A _08407_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_05596_ _05596_/A _05607_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[12\]_A3 _06840_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07335_ _07327_/CLK line[79] VGND VGND VPWR VPWR _07335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07266_ _07266_/A _07287_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_09005_ _09005_/CLK line[74] VGND VGND VPWR VPWR _09005_/Q sky130_fd_sc_hd__dfxtp_1
X_06217_ _06223_/CLK line[65] VGND VGND VPWR VPWR _06218_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07197_ _07183_/CLK line[1] VGND VGND VPWR VPWR _07197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06148_ _06147_/Q _06167_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_06079_ _06077_/CLK line[2] VGND VGND VPWR VPWR _06079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07209__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[12\].FF OVHB\[29\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[29\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09907_ _09907_/A _09912_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09838_ _09834_/CLK line[57] VGND VGND VPWR VPWR _09839_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[30\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09769_ _09768_/Q _09772_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
X_11800_ _11800_/CLK _11801_/X VGND VGND VPWR VPWR _11776_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[30\].CG clk OVHB\[30\].CGAND/X VGND VGND VPWR VPWR OVHB\[30\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_12780_ _12780_/CLK _12781_/X VGND VGND VPWR VPWR _12774_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12785__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11731_ _11872_/A wr VGND VGND VPWR VPWR _11731_/X sky130_fd_sc_hd__and2_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[15\].VALID\[7\].TOBUF OVHB\[15\].VALID\[7\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06783__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11662_ _11592_/A VGND VGND VPWR VPWR _11662_/Y sky130_fd_sc_hd__inv_2
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[23\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13400_/Q _13412_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _10627_/CLK line[32] VGND VGND VPWR VPWR _10613_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _11605_/CLK line[96] VGND VGND VPWR VPWR _11593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[2\].CG clk OVHB\[2\].CGAND/X VGND VGND VPWR VPWR OVHB\[2\].V/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10544_ _10544_/A _10577_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_13332_ _13308_/CLK line[118] VGND VGND VPWR VPWR _13332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[19\].VALID\[14\].FF OVHB\[19\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[19\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10475_ _10473_/CLK line[106] VGND VGND VPWR VPWR _10475_/Q sky130_fd_sc_hd__dfxtp_1
X_13263_ _13263_/A _13272_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_12214_ _12204_/CLK line[119] VGND VGND VPWR VPWR _12214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13194_ _13194_/CLK line[55] VGND VGND VPWR VPWR _13195_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _13900_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[22\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12025__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _12145_/A _12152_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07119__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06023__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _12072_/CLK line[56] VGND VGND VPWR VPWR _12076_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11864__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11027_ _11026_/Q _11032_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06958__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09334__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09912__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09631__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12978_ _12962_/CLK line[84] VGND VGND VPWR VPWR _12978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11929_ _11929_/A _11942_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06693__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05450_ _05449_/Q _05467_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05381_ _05391_/CLK line[67] VGND VGND VPWR VPWR _05381_/Q sky130_fd_sc_hd__dfxtp_1
X_07120_ _07120_/A _07147_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05887__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07051_ _07043_/CLK line[77] VGND VGND VPWR VPWR _07051_/Q sky130_fd_sc_hd__dfxtp_1
X_06002_ _06001_/Q _06027_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09509__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[21\].VALID\[6\].TOBUF OVHB\[21\].VALID\[6\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_115_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09806__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07953_ _07981_/CLK line[96] VGND VGND VPWR VPWR _07953_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11774__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _13515_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_56_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06904_ _06903_/Q _06937_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06868__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07884_ _07884_/A _07917_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05772__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09623_ _09622_/Q _09632_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_06835_ _06839_/CLK line[106] VGND VGND VPWR VPWR _06835_/Q sky130_fd_sc_hd__dfxtp_1
X_09554_ _09554_/CLK line[55] VGND VGND VPWR VPWR _09554_/Q sky130_fd_sc_hd__dfxtp_1
X_06766_ _06765_/Q _06797_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05717_ _05739_/CLK line[107] VGND VGND VPWR VPWR _05717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08505_ _08504_/Q _08512_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06697_ _06711_/CLK line[43] VGND VGND VPWR VPWR _06697_/Q sky130_fd_sc_hd__dfxtp_1
X_09485_ _09485_/A _09492_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07699__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08436_ _08410_/CLK line[56] VGND VGND VPWR VPWR _08436_/Q sky130_fd_sc_hd__dfxtp_1
X_05648_ _05647_/Q _05677_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[12\].FF OVHB\[1\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[1\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ _08366_/Q _08372_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XDECH.DEC0.AND2 A_h[7] A_h[8] VGND VGND VPWR VPWR _13966_/D sky130_fd_sc_hd__and2b_2
X_05579_ _05575_/CLK line[44] VGND VGND VPWR VPWR _05579_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11014__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07318_ _07292_/CLK line[57] VGND VGND VPWR VPWR _07318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06108__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08298_ _08282_/CLK line[121] VGND VGND VPWR VPWR _08298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11949__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10853__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07249_ _07248_/Q _07252_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11311__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05947__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08323__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10260_ _10260_/CLK _10261_/X VGND VGND VPWR VPWR _10248_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_105_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10191_ _10192_/A wr VGND VGND VPWR VPWR _10191_/X sky130_fd_sc_hd__and2_1
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[8\].VALID\[3\].FF OVHB\[8\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[8\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13950_ _13950_/A _13950_/B _13950_/C _13957_/D VGND VGND VPWR VPWR _13950_/Y sky130_fd_sc_hd__nor4b_4
XFILLER_4_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05682__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12901_ _12900_/Q _12922_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_13881_ _13881_/A _13902_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[17\].VALID\[12\].TOBUF OVHB\[17\].VALID\[12\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12832_ _12820_/CLK line[17] VGND VGND VPWR VPWR _12832_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _13130_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07252__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12763_ _12763_/A _12782_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11714_ _11706_/CLK line[18] VGND VGND VPWR VPWR _11715_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12708_/CLK line[82] VGND VGND VPWR VPWR _12694_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11644_/Q _11662_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11576_ _11588_/CLK line[83] VGND VGND VPWR VPWR _11576_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[25\].VALID\[10\].FF OVHB\[25\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[25\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10763__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _13314_/Q _13342_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10527_ _10527_/A _10542_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05857__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08233__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[2\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10458_ _10466_/CLK line[84] VGND VGND VPWR VPWR _10459_/A sky130_fd_sc_hd__dfxtp_1
X_13246_ _13254_/CLK line[93] VGND VGND VPWR VPWR _13246_/Q sky130_fd_sc_hd__dfxtp_1
X_13177_ _13176_/Q _13202_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_10389_ _10388_/Q _10402_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[11\].TOBUF OVHB\[10\].VALID\[11\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_124_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07427__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12128_ _12130_/CLK line[94] VGND VGND VPWR VPWR _12128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[27\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _10470_/CLK sky130_fd_sc_hd__clkbuf_4
X_12059_ _12059_/A _12082_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07146__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04950_ _04949_/Q _04977_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06688__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09064__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[20\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09999__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06620_ _06620_/CLK _06621_/X VGND VGND VPWR VPWR _06596_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10003__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06551_ _06551_/A wr VGND VGND VPWR VPWR _06551_/X sky130_fd_sc_hd__and2_1
XOVHB\[6\].VALID\[5\].FF OVHB\[6\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[6\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10938__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[12\].FF OVHB\[15\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[15\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13314__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05502_ _13908_/X VGND VGND VPWR VPWR _05502_/Y sky130_fd_sc_hd__inv_2
X_09270_ _09256_/CLK line[53] VGND VGND VPWR VPWR _09270_/Q sky130_fd_sc_hd__dfxtp_1
X_06482_ _06551_/A VGND VGND VPWR VPWR _06482_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08408__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07312__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ _08221_/A _08232_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_05433_ _05445_/CLK line[96] VGND VGND VPWR VPWR _05433_/Q sky130_fd_sc_hd__dfxtp_1
X_08152_ _08134_/CLK line[54] VGND VGND VPWR VPWR _08152_/Q sky130_fd_sc_hd__dfxtp_1
X_05364_ _05364_/A _05397_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07103_ _07103_/A _07112_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_08083_ _08082_/Q _08092_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_05295_ _05299_/CLK line[42] VGND VGND VPWR VPWR _05295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09239__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07034_ _07030_/CLK line[55] VGND VGND VPWR VPWR _07035_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08721__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13984__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08985_ _08984_/Q _09002_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06598__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07936_ _07946_/CLK line[83] VGND VGND VPWR VPWR _07937_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07867_ _07866_/Q _07882_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09606_ _09626_/CLK line[93] VGND VGND VPWR VPWR _09606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[26\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _10085_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_83_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06818_ _06802_/CLK line[84] VGND VGND VPWR VPWR _06818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07798_ _07788_/CLK line[20] VGND VGND VPWR VPWR _07798_/Q sky130_fd_sc_hd__dfxtp_1
X_09537_ _09536_/Q _09562_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_06749_ _06749_/A _06762_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _09482_/CLK line[30] VGND VGND VPWR VPWR _09468_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07222__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04938__A2_N _04938_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[23\] _13405_/Z _09555_/Z _06545_/Z _09415_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[23] sky130_fd_sc_hd__mux4_1
X_08419_ _08418_/Q _08442_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09399_ _09398_/Q _09422_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[30\].VALID\[11\].TOBUF OVHB\[30\].VALID\[11\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ _11440_/CLK line[31] VGND VGND VPWR VPWR _11430_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11679__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[7\].FF OVHB\[4\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[4\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11361_ _11361_/A _11382_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09149__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13100_ _13120_/CLK line[26] VGND VGND VPWR VPWR _13100_/Q sky130_fd_sc_hd__dfxtp_1
X_10312_ _10314_/CLK line[17] VGND VGND VPWR VPWR _10312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08053__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11976__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11292_ _11302_/CLK line[81] VGND VGND VPWR VPWR _11292_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13894__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10243_ _10242_/Q _10262_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_13031_ _13030_/Q _13062_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[25\]_A2 _13549_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[3\].TOBUF OVHB\[3\].VALID\[3\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__08988__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10174_ _10188_/CLK line[82] VGND VGND VPWR VPWR _10174_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[6\].TOBUF OVHB\[28\].VALID\[6\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12303__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06301__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13933_ _13934_/B _13933_/B _13934_/C _13934_/D VGND VGND VPWR VPWR _11032_/A sky130_fd_sc_hd__and4b_4
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VOBUF OVHB\[28\].V/Q OVHB\[28\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_13864_ _13863_/Q _13867_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10401__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09612__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12815_ _12815_/CLK _12816_/X VGND VGND VPWR VPWR _12803_/CLK sky130_fd_sc_hd__dlclkp_1
X_13795_ _13795_/CLK _13796_/X VGND VGND VPWR VPWR _13763_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_76_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12746_ _12712_/A wr VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__and2_1
XANTENNA__08228__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12712_/A VGND VGND VPWR VPWR _12677_/Y sky130_fd_sc_hd__inv_2
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _11636_/CLK line[112] VGND VGND VPWR VPWR _11628_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[15\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _06830_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10493__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11559_ _11558_/Q _11592_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05587__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[0\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05080_ _05080_/CLK _05081_/X VGND VGND VPWR VPWR _05058_/CLK sky130_fd_sc_hd__dlclkp_1
X_13229_ _13213_/CLK line[71] VGND VGND VPWR VPWR _13229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08898__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[2\].VALID\[9\].FF OVHB\[2\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[2\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06061__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05982_ _05984_/CLK line[86] VGND VGND VPWR VPWR _05982_/Q sky130_fd_sc_hd__dfxtp_1
X_08770_ _08762_/CLK line[95] VGND VGND VPWR VPWR _08770_/Q sky130_fd_sc_hd__dfxtp_1
X_04933_ A_h[21] _04933_/B2 A_h[21] _04933_/B2 VGND VGND VPWR VPWR _04936_/B sky130_fd_sc_hd__a2bb2o_4
X_07721_ _07721_/A _07742_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06211__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07652_ _07644_/CLK line[81] VGND VGND VPWR VPWR _07653_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06603_ _06602_/Q _06622_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_07583_ _07582_/Q _07602_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10668__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13044__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06534_ _06528_/CLK line[82] VGND VGND VPWR VPWR _06534_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13622__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09322_ _09320_/CLK line[91] VGND VGND VPWR VPWR _09322_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08138__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06465_ _06464_/Q _06482_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_09253_ _09253_/A _09282_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12883__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13341__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07977__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08204_ _08208_/CLK line[92] VGND VGND VPWR VPWR _08204_/Q sky130_fd_sc_hd__dfxtp_1
X_05416_ _05424_/CLK line[83] VGND VGND VPWR VPWR _05416_/Q sky130_fd_sc_hd__dfxtp_1
X_09184_ _09200_/CLK line[28] VGND VGND VPWR VPWR _09184_/Q sky130_fd_sc_hd__dfxtp_1
X_06396_ _06408_/CLK line[19] VGND VGND VPWR VPWR _06396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06236__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08135_ _08134_/Q _08162_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_05347_ _05346_/Q _05362_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_08066_ _08070_/CLK line[29] VGND VGND VPWR VPWR _08066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05278_ _05278_/CLK line[20] VGND VGND VPWR VPWR _05278_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[14\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _06445_/CLK sky130_fd_sc_hd__clkbuf_4
X_07017_ _07016_/Q _07042_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[30\].VALID\[3\].FF OVHB\[30\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[30\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08601__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13219__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[10\].FF OVHB\[11\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[11\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08968_ _08972_/CLK line[48] VGND VGND VPWR VPWR _08969_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[15\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09282__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13516__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07919_ _07918_/Q _07952_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08899_ _08898_/Q _08932_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10930_ _10930_/CLK line[58] VGND VGND VPWR VPWR _10930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05960__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10578__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10861_ _10861_/A _10892_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_12600_ _12599_/Q _12607_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[8\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13580_ _13580_/A _13587_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[27\].CGAND_A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10792_ _10804_/CLK line[123] VGND VGND VPWR VPWR _10792_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[8\].TOBUF OVHB\[1\].VALID\[8\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12531_ _12523_/CLK line[8] VGND VGND VPWR VPWR _12531_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12793__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07887__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06791__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12462_ _12462_/A _12467_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11413_ _11395_/CLK line[9] VGND VGND VPWR VPWR _11413_/Q sky130_fd_sc_hd__dfxtp_1
X_12393_ _12387_/CLK line[73] VGND VGND VPWR VPWR _12393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10891__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09457__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11344_ _11344_/A _11347_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[4\].FF OVHB\[29\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[29\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05200__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09176__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11275_ _11275_/CLK _11276_/X VGND VGND VPWR VPWR _11251_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_79_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13014_ _13013_/Q _13027_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10226_ _10192_/A wr VGND VGND VPWR VPWR _10226_/X sky130_fd_sc_hd__and2_1
XANTENNA__12033__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10157_ _10192_/A VGND VGND VPWR VPWR _10157_/Y sky130_fd_sc_hd__inv_2
XOVHB\[11\].VALID\[1\].FF OVHB\[11\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[11\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07127__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10088_ _10100_/CLK line[48] VGND VGND VPWR VPWR _10088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12968__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06966__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13916_ A[6] VGND VGND VPWR VPWR _13923_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__09342__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13847_ _13845_/CLK line[97] VGND VGND VPWR VPWR _13847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[17\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13778_ _13777_/Q _13797_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_12729_ _12741_/CLK line[98] VGND VGND VPWR VPWR _12729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06250_ _06244_/CLK line[95] VGND VGND VPWR VPWR _06250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05201_ _05200_/Q _05222_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
X_06181_ _06180_/Q _06202_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12208__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04940__A1_N A_h[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05132_ _05122_/CLK line[81] VGND VGND VPWR VPWR _05132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09940_ _09939_/Q _09947_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_05063_ _05063_/A _05082_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09517__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09871_ _09849_/CLK line[72] VGND VGND VPWR VPWR _09871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[28\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08822_ _08821_/Q _08827_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[6\].FF OVHB\[27\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[27\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[14\].TOBUF OVHB\[7\].VALID\[14\].FF/Q OVHB\[7\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_08753_ _08749_/CLK line[73] VGND VGND VPWR VPWR _08754_/A sky130_fd_sc_hd__dfxtp_1
X_05965_ _05965_/A _05992_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11782__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07704_ _07703_/Q _07707_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11137__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04916_ _04915_/Y _04918_/B2 _04916_/B1 VGND VGND VPWR VPWR _04916_/X sky130_fd_sc_hd__o21a_4
XOVHB\[6\].VALID\[12\].FF OVHB\[6\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[6\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[7\]_A2 _13510_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06876__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08684_ _08683_/Q _08687_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_05896_ _05902_/CLK line[61] VGND VGND VPWR VPWR _05896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09252__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10398__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07635_ _07635_/CLK _07636_/X VGND VGND VPWR VPWR _07633_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[15\]_A1 _05586_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07566_ _07672_/A wr VGND VGND VPWR VPWR _07566_/X sky130_fd_sc_hd__and2_1
XFILLER_0_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09305_ _09307_/CLK line[69] VGND VGND VPWR VPWR _09305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06517_ _06551_/A VGND VGND VPWR VPWR _06517_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07497_ _07672_/A VGND VGND VPWR VPWR _07497_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09236_ _09235_/Q _09247_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_06448_ _06464_/CLK line[48] VGND VGND VPWR VPWR _06449_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07500__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12118__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09167_ _09147_/CLK line[6] VGND VGND VPWR VPWR _09168_/A sky130_fd_sc_hd__dfxtp_1
X_06379_ _06378_/Q _06412_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11022__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08118_ _08117_/Q _08127_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06116__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09098_ _09098_/A _09107_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[10\].TOBUF OVHB\[27\].VALID\[10\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11957__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[13\].TOBUF OVHB\[0\].VALID\[13\].FF/Q OVHB\[0\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08049_ _08033_/CLK line[7] VGND VGND VPWR VPWR _08049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09427__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11060_ _11060_/A _11067_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08331__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10011_ _10011_/CLK line[8] VGND VGND VPWR VPWR _10011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12431__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11962_ _11961_/Q _11977_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05690__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13701_ _13701_/CLK line[45] VGND VGND VPWR VPWR _13702_/A sky130_fd_sc_hd__dfxtp_1
X_10913_ _10903_/CLK line[36] VGND VGND VPWR VPWR _10913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11893_ _11901_/CLK line[100] VGND VGND VPWR VPWR _11894_/A sky130_fd_sc_hd__dfxtp_1
X_13632_ _13632_/A _13657_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[8\].FF OVHB\[25\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[25\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10844_ _10844_/A _10857_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_13563_ _13559_/CLK line[110] VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__dfxtp_1
X_10775_ _10783_/CLK line[101] VGND VGND VPWR VPWR _10775_/Q sky130_fd_sc_hd__dfxtp_1
X_12514_ _12513_/Q _12537_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08506__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13494_ _13493_/Q _13517_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ _12449_/CLK line[111] VGND VGND VPWR VPWR _12445_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12606__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ _12375_/Q _12397_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08091__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10771__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11327_ _11343_/CLK line[97] VGND VGND VPWR VPWR _11327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05865__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08241__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11258_ _11257_/Q _11277_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_10209_ _10217_/CLK line[98] VGND VGND VPWR VPWR _10210_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11189_ _11191_/CLK line[34] VGND VGND VPWR VPWR _11189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12698__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05750_ _05756_/CLK line[122] VGND VGND VPWR VPWR _05750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05681_ _05681_/A _05712_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11107__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07420_ _07419_/Q _07427_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10011__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08266__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05105__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10946__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07351_ _07327_/CLK line[72] VGND VGND VPWR VPWR _07351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13322__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06302_ _06301_/Q _06307_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
X_07282_ _07281_/Q _07287_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08416__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[8\].TOBUF OVHB\[8\].VALID\[8\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_06233_ _06223_/CLK line[73] VGND VGND VPWR VPWR _06233_/Q sky130_fd_sc_hd__dfxtp_1
X_09021_ _09005_/CLK line[67] VGND VGND VPWR VPWR _09022_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06164_ _06163_/Q _06167_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_05115_ _05115_/CLK _05116_/X VGND VGND VPWR VPWR _05093_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06095_ _06095_/CLK _06096_/X VGND VGND VPWR VPWR _06077_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_132_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09923_ _09925_/CLK line[110] VGND VGND VPWR VPWR _09924_/A sky130_fd_sc_hd__dfxtp_1
X_05046_ _05152_/A wr VGND VGND VPWR VPWR _05046_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[11\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09854_ _09854_/A _09877_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07990__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08805_ _08823_/CLK line[111] VGND VGND VPWR VPWR _08805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09785_ _09793_/CLK line[47] VGND VGND VPWR VPWR _09785_/Q sky130_fd_sc_hd__dfxtp_1
X_06997_ _07001_/CLK line[38] VGND VGND VPWR VPWR _06997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08736_ _08735_/Q _08757_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05948_ _05948_/A _05957_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08667_ _08663_/CLK line[33] VGND VGND VPWR VPWR _08667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05879_ _05871_/CLK line[39] VGND VGND VPWR VPWR _05879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07618_ _07617_/Q _07637_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05015__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08598_ _08597_/Q _08617_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _07539_/CLK line[34] VGND VGND VPWR VPWR _07549_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560_ _10559_/Q _10577_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07230__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[30\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09219_ _09241_/CLK line[44] VGND VGND VPWR VPWR _09219_/Q sky130_fd_sc_hd__dfxtp_1
X_10491_ _10473_/CLK line[99] VGND VGND VPWR VPWR _10491_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _12745_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_33_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ _12229_/Q _12257_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11687__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12161_ _12177_/CLK line[109] VGND VGND VPWR VPWR _12161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[10\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09157__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11112_ _11112_/A _11137_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[10\].FF OVHB\[2\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[2\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12092_ _12092_/A _12117_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[3\].TOBUF OVHB\[15\].VALID\[3\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08996__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11043_ _11063_/CLK line[110] VGND VGND VPWR VPWR _11043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12311__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12994_ _12993_/Q _13027_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07405__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DEC.DEC0.AND1_B A[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11945_ _11945_/CLK line[10] VGND VGND VPWR VPWR _11946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11876_ _11876_/A _11907_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09620__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13615_ _13615_/A _13622_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_10827_ _10843_/CLK line[11] VGND VGND VPWR VPWR _10827_/Q sky130_fd_sc_hd__dfxtp_1
X_13546_ _13528_/CLK line[88] VGND VGND VPWR VPWR _13546_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10758_ _10757_/Q _10787_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_13477_ _13476_/Q _13482_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_10689_ _10707_/CLK line[76] VGND VGND VPWR VPWR _10689_/Q sky130_fd_sc_hd__dfxtp_1
X_12428_ _12414_/CLK line[89] VGND VGND VPWR VPWR _12428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11597__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12359_ _12359_/A _12362_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05595__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[4\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _12360_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_49_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13167__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06920_ _06920_/A _06937_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06851_ _06839_/CLK line[99] VGND VGND VPWR VPWR _06851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05802_ _05801_/Q _05817_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09570_ _09570_/A _09597_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_06782_ _06782_/A _06797_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_08521_ _08541_/CLK line[109] VGND VGND VPWR VPWR _08521_/Q sky130_fd_sc_hd__dfxtp_1
X_05733_ _05739_/CLK line[100] VGND VGND VPWR VPWR _05734_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[2\].TOBUF OVHB\[21\].VALID\[2\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_08452_ _08451_/Q _08477_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
X_05664_ _05663_/Q _05677_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09530__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07403_ _07393_/CLK line[110] VGND VGND VPWR VPWR _07404_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10676__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[20\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08383_ _08383_/CLK line[46] VGND VGND VPWR VPWR _08384_/A sky130_fd_sc_hd__dfxtp_1
X_05595_ _05575_/CLK line[37] VGND VGND VPWR VPWR _05596_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13052__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[29\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08146__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07334_ _07333_/Q _07357_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13987__D _13990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07265_ _07267_/CLK line[47] VGND VGND VPWR VPWR _07266_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _09700_/CLK sky130_fd_sc_hd__clkbuf_4
X_09004_ _09003_/Q _09037_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_06216_ _06216_/A _06237_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_07196_ _07195_/Q _07217_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[29\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[10\].FF OVHB\[16\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[16\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06147_ _06147_/CLK line[33] VGND VGND VPWR VPWR _06147_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11300__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06078_ _06077_/Q _06097_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05029_ _05041_/CLK line[34] VGND VGND VPWR VPWR _05029_/Q sky130_fd_sc_hd__dfxtp_1
X_09906_ _09908_/CLK line[88] VGND VGND VPWR VPWR _09907_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09705__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09837_ _09837_/A _09842_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDATA\[3\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _11975_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13227__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09768_ _09760_/CLK line[25] VGND VGND VPWR VPWR _09768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08719_ _08718_/Q _08722_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_09699_ _09699_/A _09702_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11730_ _11730_/CLK _11731_/X VGND VGND VPWR VPWR _11706_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10586__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _11592_/A wr VGND VGND VPWR VPWR _11661_/X sky130_fd_sc_hd__and2_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13394_/CLK line[21] VGND VGND VPWR VPWR _13400_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[8\].TOBUF OVHB\[13\].VALID\[8\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_10612_ _13932_/X VGND VGND VPWR VPWR _10612_/Y sky130_fd_sc_hd__inv_2
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _11592_/A VGND VGND VPWR VPWR _11592_/Y sky130_fd_sc_hd__inv_2
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13331_ _13330_/Q _13342_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_10543_ _10571_/CLK line[0] VGND VGND VPWR VPWR _10544_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13262_ _13254_/CLK line[86] VGND VGND VPWR VPWR _13263_/A sky130_fd_sc_hd__dfxtp_1
X_10474_ _10474_/A _10507_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[28\]_A0 _10865_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12213_ _12212_/Q _12222_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_13193_ _13192_/Q _13202_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11210__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[23\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _09315_/CLK sky130_fd_sc_hd__clkbuf_4
X_12144_ _12130_/CLK line[87] VGND VGND VPWR VPWR _12145_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12075_ _12075_/A _12082_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_11026_ _11002_/CLK line[88] VGND VGND VPWR VPWR _11026_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13137__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12041__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07135__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12976__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12977_ _12977_/A _12992_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11928_ _11934_/CLK line[116] VGND VGND VPWR VPWR _11929_/A sky130_fd_sc_hd__dfxtp_1
X_11859_ _11858_/Q _11872_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05380_ _05379_/Q _05397_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13529_ _13528_/Q _13552_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13600__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07050_ _07049_/Q _07077_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06001_ _06023_/CLK line[109] VGND VGND VPWR VPWR _06001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12216__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07952_ _13920_/X VGND VGND VPWR VPWR _07952_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[17\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06903_ _06923_/CLK line[0] VGND VGND VPWR VPWR _06903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07883_ _07905_/CLK line[64] VGND VGND VPWR VPWR _07884_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _08930_/CLK sky130_fd_sc_hd__clkbuf_4
X_09622_ _09626_/CLK line[86] VGND VGND VPWR VPWR _09622_/Q sky130_fd_sc_hd__dfxtp_1
X_06834_ _06833_/Q _06867_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07045__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09553_ _09553_/A _09562_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[12\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _06060_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_71_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06765_ _06775_/CLK line[74] VGND VGND VPWR VPWR _06765_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11790__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08504_ _08480_/CLK line[87] VGND VGND VPWR VPWR _08504_/Q sky130_fd_sc_hd__dfxtp_1
X_05716_ _05716_/A _05747_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06884__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _09482_/CLK line[23] VGND VGND VPWR VPWR _09485_/A sky130_fd_sc_hd__dfxtp_1
X_06696_ _06696_/A _06727_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09260__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08435_ _08434_/Q _08442_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_05647_ _05671_/CLK line[75] VGND VGND VPWR VPWR _05647_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[27\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ _08358_/CLK line[24] VGND VGND VPWR VPWR _08366_/Q sky130_fd_sc_hd__dfxtp_1
X_05578_ _05577_/Q _05607_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XDECH.DEC0.AND3 A_h[8] A_h[7] VGND VGND VPWR VPWR _13979_/D sky130_fd_sc_hd__and2_2
X_07317_ _07316_/Q _07322_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08297_ _08296_/Q _08302_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_07248_ _07232_/CLK line[25] VGND VGND VPWR VPWR _07248_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12126__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07179_ _07178_/Q _07182_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06124__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10190_ _10190_/CLK _10191_/X VGND VGND VPWR VPWR _10188_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11965__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[13\].TOBUF OVHB\[13\].VALID\[13\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09435__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _12902_/CLK line[63] VGND VGND VPWR VPWR _12900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13880_ _13882_/CLK line[127] VGND VGND VPWR VPWR _13881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12831_ _12830_/Q _12852_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12762_ _12774_/CLK line[113] VGND VGND VPWR VPWR _12763_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11712_/Q _11732_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12692_/Q _12712_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[11\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _05675_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[2\].TOBUF OVHB\[28\].VALID\[2\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11636_/CLK line[114] VGND VGND VPWR VPWR _11644_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[18\].INV _13963_/X VGND VGND VPWR VPWR OVHB\[18\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11574_/Q _11592_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13314_ _13308_/CLK line[124] VGND VGND VPWR VPWR _13314_/Q sky130_fd_sc_hd__dfxtp_1
X_10526_ _10520_/CLK line[115] VGND VGND VPWR VPWR _10527_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VOBUF OVHB\[24\].V/Q OVHB\[24\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13245_ _13244_/Q _13272_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[2\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10457_ _10456_/Q _10472_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06034__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13176_ _13194_/CLK line[61] VGND VGND VPWR VPWR _13176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10388_ _10384_/CLK line[52] VGND VGND VPWR VPWR _10388_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11875__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[0\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12127_ _12127_/A _12152_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[10\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05873__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12058_ _12072_/CLK line[62] VGND VGND VPWR VPWR _12059_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11009_ _11008_/Q _11032_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06550_ _06550_/CLK _06551_/X VGND VGND VPWR VPWR _06528_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_34_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05501_ _13908_/X wr VGND VGND VPWR VPWR _05501_/X sky130_fd_sc_hd__and2_1
X_06481_ _06551_/A wr VGND VGND VPWR VPWR _06481_/X sky130_fd_sc_hd__and2_1
XANTENNA__11115__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08220_ _08208_/CLK line[85] VGND VGND VPWR VPWR _08221_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06209__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05432_ _13908_/X VGND VGND VPWR VPWR _05432_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05113__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08151_ _08150_/Q _08162_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10954__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05363_ _05391_/CLK line[64] VGND VGND VPWR VPWR _05364_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13330__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07102_ _07098_/CLK line[86] VGND VGND VPWR VPWR _07103_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08424__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _05290_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05294_ _05293_/Q _05327_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_08082_ _08070_/CLK line[22] VGND VGND VPWR VPWR _08082_/Q sky130_fd_sc_hd__dfxtp_1
X_07033_ _07032_/Q _07042_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08721__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].CG clk OVHB\[20\].CG/GATE VGND VGND VPWR VPWR OVHB\[20\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_115_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ _08972_/CLK line[50] VGND VGND VPWR VPWR _08984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05783__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07935_ _07934_/Q _07952_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[1\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07866_ _07854_/CLK line[51] VGND VGND VPWR VPWR _07866_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04977__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09605_ _09604_/Q _09632_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06817_ _06816_/Q _06832_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07797_ _07796_/Q _07812_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13505__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09536_ _09554_/CLK line[61] VGND VGND VPWR VPWR _09536_/Q sky130_fd_sc_hd__dfxtp_1
X_06748_ _06740_/CLK line[52] VGND VGND VPWR VPWR _06749_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ _09466_/Q _09492_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_06679_ _06679_/A _06692_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ _08410_/CLK line[62] VGND VGND VPWR VPWR _08418_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05023__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09398_ _09414_/CLK line[126] VGND VGND VPWR VPWR _09398_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10864__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ _08348_/Q _08372_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[16\] _10859_/Z _07009_/Z _05119_/Z _13589_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[16] sky130_fd_sc_hd__mux4_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05958__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13240__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[10\].FF OVHB\[7\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[7\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11360_ _11370_/CLK line[127] VGND VGND VPWR VPWR _11361_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10311_ _10310_/Q _10332_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11291_ _11290_/Q _11312_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13030_ _13050_/CLK line[122] VGND VGND VPWR VPWR _13030_/Q sky130_fd_sc_hd__dfxtp_1
X_10242_ _10248_/CLK line[113] VGND VGND VPWR VPWR _10242_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[25\]_A3 _07179_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[1\].VALID\[4\].TOBUF OVHB\[1\].VALID\[4\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06789__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10173_ _10173_/A _10192_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09165__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[7\].TOBUF OVHB\[26\].VALID\[7\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_121_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[25\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10104__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13932_ _13933_/B _13934_/B _13934_/C _13934_/D VGND VGND VPWR VPWR _13932_/X sky130_fd_sc_hd__and4bb_4
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13863_ _13845_/CLK line[105] VGND VGND VPWR VPWR _13863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13415__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10401__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _12814_/A _12817_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_13794_ _13793_/Q _13797_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07413__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12745_ _12745_/CLK _12746_/X VGND VGND VPWR VPWR _12741_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_70_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12712_/A wr VGND VGND VPWR VPWR _12676_/X sky130_fd_sc_hd__and2_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _11592_/A VGND VGND VPWR VPWR _11627_/Y sky130_fd_sc_hd__inv_2
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _11588_/CLK line[80] VGND VGND VPWR VPWR _11558_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[2\].FF OVHB\[18\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[18\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10509_ _10508_/Q _10542_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
X_11489_ _11488_/Q _11522_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_13228_ _13227_/Q _13237_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06342__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13159_ _13163_/CLK line[39] VGND VGND VPWR VPWR _13159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06699__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09075__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06061__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05981_ _05981_/A _05992_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_07720_ _07724_/CLK line[127] VGND VGND VPWR VPWR _07721_/A sky130_fd_sc_hd__dfxtp_1
X_04932_ A_h[11] _04932_/B2 A_h[11] _04932_/B2 VGND VGND VPWR VPWR _04932_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__09803__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07651_ _07650_/Q _07672_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06602_ _06596_/CLK line[113] VGND VGND VPWR VPWR _06602_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04947__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13903__A A[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07582_ _07572_/CLK line[49] VGND VGND VPWR VPWR _07582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07323__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09321_ _09320_/Q _09352_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_06533_ _06532_/Q _06552_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09252_ _09256_/CLK line[59] VGND VGND VPWR VPWR _09253_/A sky130_fd_sc_hd__dfxtp_1
X_06464_ _06464_/CLK line[50] VGND VGND VPWR VPWR _06464_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06517__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08203_ _08202_/Q _08232_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_05415_ _05414_/Q _05432_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_09183_ _09182_/Q _09212_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_06395_ _06395_/A _06412_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06236__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05778__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[10\].TOBUF OVHB\[7\].VALID\[10\].FF/Q OVHB\[7\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_08134_ _08134_/CLK line[60] VGND VGND VPWR VPWR _08134_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08154__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05346_ _05332_/CLK line[51] VGND VGND VPWR VPWR _05346_/Q sky130_fd_sc_hd__dfxtp_1
X_08065_ _08064_/Q _08092_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_05277_ _05276_/Q _05292_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_07016_ _07030_/CLK line[61] VGND VGND VPWR VPWR _07016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12404__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[16\].VALID\[4\].FF OVHB\[16\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[16\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06402__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08967_ _13923_/X VGND VGND VPWR VPWR _08967_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07918_ _07946_/CLK line[80] VGND VGND VPWR VPWR _07918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08898_ _08922_/CLK line[16] VGND VGND VPWR VPWR _08898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09713__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07849_ _07848_/Q _07882_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08329__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10860_ _10872_/CLK line[26] VGND VGND VPWR VPWR _10861_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ _09507_/CLK line[39] VGND VGND VPWR VPWR _09520_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07811__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10791_ _10790_/Q _10822_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[27\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12529_/Q _12537_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10594__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12461_ _12449_/CLK line[104] VGND VGND VPWR VPWR _12462_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05688__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11412_ _11411_/Q _11417_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08064__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12392_ _12391_/Q _12397_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10891__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11343_ _11343_/CLK line[105] VGND VGND VPWR VPWR _11344_/A sky130_fd_sc_hd__dfxtp_1
X_11274_ _11273_/Q _11277_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_13013_ _12999_/CLK line[100] VGND VGND VPWR VPWR _13013_/Q sky130_fd_sc_hd__dfxtp_1
X_10225_ _10225_/CLK _10226_/X VGND VGND VPWR VPWR _10217_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06312__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10156_ _10192_/A wr VGND VGND VPWR VPWR _10156_/X sky130_fd_sc_hd__and2_1
X_10087_ _10192_/A VGND VGND VPWR VPWR _10087_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[29\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10769__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13915_ A[5] VGND VGND VPWR VPWR _13923_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13145__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08239__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13846_ _13846_/A _13867_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[6\].FF OVHB\[14\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[14\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07143__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12984__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[23\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13777_ _13763_/CLK line[65] VGND VGND VPWR VPWR _13777_/Q sky130_fd_sc_hd__dfxtp_1
X_10989_ _10977_/CLK line[71] VGND VGND VPWR VPWR _10989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12728_ _12727_/Q _12747_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _12667_/CLK line[66] VGND VGND VPWR VPWR _12659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05200_ _05214_/CLK line[127] VGND VGND VPWR VPWR _05200_/Q sky130_fd_sc_hd__dfxtp_1
X_06180_ _06186_/CLK line[63] VGND VGND VPWR VPWR _06180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05131_ _05130_/Q _05152_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10009__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05062_ _05058_/CLK line[49] VGND VGND VPWR VPWR _05063_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08702__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09870_ _09869_/Q _09877_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07318__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08821_ _08823_/CLK line[104] VGND VGND VPWR VPWR _08821_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04937__A2_N _04937_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[8\].VALID\[4\].TOBUF OVHB\[8\].VALID\[4\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_135_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08752_ _08752_/A _08757_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_05964_ _05984_/CLK line[92] VGND VGND VPWR VPWR _05965_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07703_ _07679_/CLK line[105] VGND VGND VPWR VPWR _07703_/Q sky130_fd_sc_hd__dfxtp_1
X_04915_ A_h[18] VGND VGND VPWR VPWR _04915_/Y sky130_fd_sc_hd__inv_2
X_08683_ _08663_/CLK line[41] VGND VGND VPWR VPWR _08683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[7\]_A3 _07140_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05895_ _05894_/Q _05922_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07634_ _07633_/Q _07637_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07053__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12894__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07565_ _07565_/CLK _07566_/X VGND VGND VPWR VPWR _07539_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.MUX\[15\]_A2 _13496_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07988__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09304_ _09303_/Q _09317_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_06516_ _06551_/A wr VGND VGND VPWR VPWR _06516_/X sky130_fd_sc_hd__and2_1
XANTENNA__06892__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07496_ _07672_/A wr VGND VGND VPWR VPWR _07496_/X sky130_fd_sc_hd__and2_1
XOVHB\[23\].VALID\[11\].TOBUF OVHB\[23\].VALID\[11\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05151__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09235_ _09241_/CLK line[37] VGND VGND VPWR VPWR _09235_/Q sky130_fd_sc_hd__dfxtp_1
X_06447_ _06551_/A VGND VGND VPWR VPWR _06447_/Y sky130_fd_sc_hd__inv_2
XDATA\[1\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _08230_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[12\].VALID\[8\].FF OVHB\[12\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[12\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09166_ _09165_/Q _09177_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_06378_ _06408_/CLK line[16] VGND VGND VPWR VPWR _06378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05301__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08117_ _08113_/CLK line[38] VGND VGND VPWR VPWR _08117_/Q sky130_fd_sc_hd__dfxtp_1
X_05329_ _05328_/Q _05362_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09097_ _09085_/CLK line[102] VGND VGND VPWR VPWR _09098_/A sky130_fd_sc_hd__dfxtp_1
X_08048_ _08047_/Q _08057_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12134__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12712__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07228__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10010_ _10009_/Q _10017_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09999_ _10011_/CLK line[2] VGND VGND VPWR VPWR _10000_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11973__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12431__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09443__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[31\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _11800_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05326__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11961_ _11945_/CLK line[3] VGND VGND VPWR VPWR _11961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ _13699_/Q _13727_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_10912_ _10911_/Q _10927_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11892_ _11891_/Q _11907_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
X_13631_ _13631_/CLK line[13] VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10843_ _10843_/CLK line[4] VGND VGND VPWR VPWR _10844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13562_ _13561_/Q _13587_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_10774_ _10773_/Q _10787_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
X_12513_ _12523_/CLK line[14] VGND VGND VPWR VPWR _12513_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12309__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13493_ _13497_/CLK line[78] VGND VGND VPWR VPWR _13493_/Q sky130_fd_sc_hd__dfxtp_1
X_12444_ _12443_/Q _12467_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08372__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12606__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _12387_/CLK line[79] VGND VGND VPWR VPWR _12375_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[0\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _05045_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08091__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09618__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11326_ _11326_/A _11347_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11257_ _11251_/CLK line[65] VGND VGND VPWR VPWR _11257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[25\].V OVHB\[25\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[25\].V/Q sky130_fd_sc_hd__dfrtp_1
X_10208_ _10208_/A _10227_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06042__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11188_ _11188_/A _11207_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11883__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06977__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10139_ _10145_/CLK line[66] VGND VGND VPWR VPWR _10139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05881__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09353__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[3\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10499__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05680_ _05708_/CLK line[90] VGND VGND VPWR VPWR _05681_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08547__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13829_ _13829_/A _13832_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08266__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _11415_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07350_ _07349_/Q _07357_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_06301_ _06285_/CLK line[104] VGND VGND VPWR VPWR _06301_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[20\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _08545_/CLK sky130_fd_sc_hd__clkbuf_4
X_07281_ _07267_/CLK line[40] VGND VGND VPWR VPWR _07281_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11123__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09020_ _09019_/Q _09037_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_06232_ _06231_/Q _06237_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[9\].TOBUF OVHB\[6\].VALID\[9\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06217__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06163_ _06147_/CLK line[41] VGND VGND VPWR VPWR _06163_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09528__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05114_ _05113_/Q _05117_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08432__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06094_ _06093_/Q _06097_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09922_ _09921_/Q _09947_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
X_05045_ _05045_/CLK _05046_/X VGND VGND VPWR VPWR _05041_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[16\].V OVHB\[16\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[16\].V/Q sky130_fd_sc_hd__dfrtp_1
X_09853_ _09849_/CLK line[78] VGND VGND VPWR VPWR _09854_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08804_ _08803_/Q _08827_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_09784_ _09783_/Q _09807_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10052__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04918__B2 _04918_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06996_ _06995_/Q _07007_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05791__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09841__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08735_ _08749_/CLK line[79] VGND VGND VPWR VPWR _08735_/Q sky130_fd_sc_hd__dfxtp_1
X_05947_ _05929_/CLK line[70] VGND VGND VPWR VPWR _05948_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[25\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08666_ _08665_/Q _08687_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_05878_ _05877_/Q _05887_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
X_07617_ _07633_/CLK line[65] VGND VGND VPWR VPWR _07617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08597_ _08609_/CLK line[1] VGND VGND VPWR VPWR _08597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13513__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _07548_/A _07567_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08607__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[18\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07479_ _07467_/CLK line[2] VGND VGND VPWR VPWR _07479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11033__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09218_ _09217_/Q _09247_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_10490_ _10489_/Q _10507_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05031__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[1\].FF OVHB\[5\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[5\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09149_ _09147_/CLK line[12] VGND VGND VPWR VPWR _09149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10872__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10227__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05966__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12160_ _12159_/Q _12187_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08342__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11111_ _11111_/CLK line[13] VGND VGND VPWR VPWR _11112_/A sky130_fd_sc_hd__dfxtp_1
X_12091_ _12109_/CLK line[77] VGND VGND VPWR VPWR _12092_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11042_ _11041_/Q _11067_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12799__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[13\].VALID\[4\].TOBUF OVHB\[13\].VALID\[4\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09173__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11208__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12993_ _12999_/CLK line[96] VGND VGND VPWR VPWR _12993_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10112__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11944_ _11943_/Q _11977_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05206__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11875_ _11901_/CLK line[106] VGND VGND VPWR VPWR _11876_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13423__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10826_ _10825_/Q _10857_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_13614_ _13598_/CLK line[119] VGND VGND VPWR VPWR _13615_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08517__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07421__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12039__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13545_ _13544_/Q _13552_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_10757_ _10783_/CLK line[107] VGND VGND VPWR VPWR _10757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11521__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13476_ _13468_/CLK line[56] VGND VGND VPWR VPWR _13476_/Q sky130_fd_sc_hd__dfxtp_1
X_10688_ _10687_/Q _10717_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12427_ _12427_/A _12432_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[16\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09348__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12358_ _12352_/CLK line[57] VGND VGND VPWR VPWR _12359_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11309_ _11309_/A _11312_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_12289_ _12288_/Q _12292_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[3\].VALID\[3\].FF OVHB\[3\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[3\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06850_ _06850_/A _06867_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09083__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05801_ _05799_/CLK line[3] VGND VGND VPWR VPWR _05801_/Q sky130_fd_sc_hd__dfxtp_1
X_06781_ _06775_/CLK line[67] VGND VGND VPWR VPWR _06782_/A sky130_fd_sc_hd__dfxtp_1
X_08520_ _08519_/Q _08547_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10022__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].VOBUF OVHB\[19\].V/Q OVHB\[19\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_05732_ _05731_/Q _05747_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07181__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08451_ _08473_/CLK line[77] VGND VGND VPWR VPWR _08451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05663_ _05671_/CLK line[68] VGND VGND VPWR VPWR _05663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07402_ _07401_/Q _07427_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04955__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08382_ _08381_/Q _08407_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_05594_ _05593_/Q _05607_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07331__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07333_ _07327_/CLK line[78] VGND VGND VPWR VPWR _07333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ _07263_/Q _07287_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11788__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09003_ _09005_/CLK line[64] VGND VGND VPWR VPWR _09003_/Q sky130_fd_sc_hd__dfxtp_1
X_06215_ _06223_/CLK line[79] VGND VGND VPWR VPWR _06216_/A sky130_fd_sc_hd__dfxtp_1
X_07195_ _07183_/CLK line[15] VGND VGND VPWR VPWR _07195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09258__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06146_ _06146_/A _06167_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06077_ _06077_/CLK line[1] VGND VGND VPWR VPWR _06077_/Q sky130_fd_sc_hd__dfxtp_1
X_05028_ _05027_/Q _05047_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07356__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09905_ _09904_/Q _09912_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12412__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09836_ _09834_/CLK line[56] VGND VGND VPWR VPWR _09837_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07506__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06979_ _07001_/CLK line[44] VGND VGND VPWR VPWR _06979_/Q sky130_fd_sc_hd__dfxtp_1
X_09767_ _09766_/Q _09772_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11028__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08718_ _08710_/CLK line[57] VGND VGND VPWR VPWR _08718_/Q sky130_fd_sc_hd__dfxtp_1
X_09698_ _09694_/CLK line[121] VGND VGND VPWR VPWR _09699_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09721__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[1\].VALID\[5\].FF OVHB\[1\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[1\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08649_ _08648_/Q _08652_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _11660_/CLK _11661_/X VGND VGND VPWR VPWR _11636_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _13932_/X wr VGND VGND VPWR VPWR _10611_/X sky130_fd_sc_hd__and2_1
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _11592_/A wr VGND VGND VPWR VPWR _11591_/X sky130_fd_sc_hd__and2_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[11\].VALID\[9\].TOBUF OVHB\[11\].VALID\[9\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_13330_ _13308_/CLK line[117] VGND VGND VPWR VPWR _13330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ _13931_/X VGND VGND VPWR VPWR _10542_/Y sky130_fd_sc_hd__inv_2
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11698__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13260_/Q _13272_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10473_ _10473_/CLK line[96] VGND VGND VPWR VPWR _10474_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05696__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12212_ _12204_/CLK line[118] VGND VGND VPWR VPWR _12212_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[28\]_A1 _07015_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08072__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13192_ _13194_/CLK line[54] VGND VGND VPWR VPWR _13192_/Q sky130_fd_sc_hd__dfxtp_1
X_12143_ _12142_/Q _12152_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12074_ _12072_/CLK line[55] VGND VGND VPWR VPWR _12075_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11025_ _11025_/A _11032_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06320__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[20\].VOBUF OVHB\[20\].V/Q OVHB\[20\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_12976_ _12962_/CLK line[83] VGND VGND VPWR VPWR _12977_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10777__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11927_ _11927_/A _11942_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13153__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08247__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11858_ _11846_/CLK line[84] VGND VGND VPWR VPWR _11858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10809_ _10808_/Q _10822_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_11789_ _11788_/Q _11802_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ _13528_/CLK line[94] VGND VGND VPWR VPWR _13528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13459_ _13458_/Q _13482_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11401__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06000_ _06000_/A _06027_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12082__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08710__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07951_ _13920_/X wr VGND VGND VPWR VPWR _07951_/X sky130_fd_sc_hd__and2_1
XANTENNA__13328__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[14\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06902_ _06832_/A VGND VGND VPWR VPWR _06902_/Y sky130_fd_sc_hd__inv_2
X_07882_ _13920_/X VGND VGND VPWR VPWR _07882_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[21\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[0\].FF OVHB\[28\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[28\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06833_ _06839_/CLK line[96] VGND VGND VPWR VPWR _06833_/Q sky130_fd_sc_hd__dfxtp_1
X_09621_ _09621_/A _09632_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09552_ _09554_/CLK line[54] VGND VGND VPWR VPWR _09553_/A sky130_fd_sc_hd__dfxtp_1
X_06764_ _06763_/Q _06797_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08503_ _08503_/A _08512_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_05715_ _05739_/CLK line[106] VGND VGND VPWR VPWR _05716_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10687__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09483_ _09482_/Q _09492_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_06695_ _06711_/CLK line[42] VGND VGND VPWR VPWR _06696_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13063__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08434_ _08410_/CLK line[55] VGND VGND VPWR VPWR _08434_/Q sky130_fd_sc_hd__dfxtp_1
X_05646_ _05645_/Q _05677_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07061__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ _08364_/Q _08372_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_05577_ _05575_/CLK line[43] VGND VGND VPWR VPWR _05577_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07996__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07316_ _07292_/CLK line[56] VGND VGND VPWR VPWR _07316_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[7\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08296_ _08282_/CLK line[120] VGND VGND VPWR VPWR _08296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ _07246_/Q _07252_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _07170_/CLK line[121] VGND VGND VPWR VPWR _07178_/Q sky130_fd_sc_hd__dfxtp_1
X_06129_ _06128_/Q _06132_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08620__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13238__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12142__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07236__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[19\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09819_ _09819_/A _09842_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12830_ _12820_/CLK line[31] VGND VGND VPWR VPWR _12830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09451__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12760_/Q _12782_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13551__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11706_/CLK line[17] VGND VGND VPWR VPWR _11712_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12708_/CLK line[81] VGND VGND VPWR VPWR _12692_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[21\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[0\].TOBUF OVHB\[1\].VALID\[0\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[2\].FF OVHB\[26\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[26\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A _11662_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[2\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13701__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[26\].VALID\[3\].TOBUF OVHB\[26\].VALID\[3\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _11588_/CLK line[82] VGND VGND VPWR VPWR _11574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13313_/A _13342_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
X_10525_ _10524_/Q _10542_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12317__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13244_ _13254_/CLK line[92] VGND VGND VPWR VPWR _13244_/Q sky130_fd_sc_hd__dfxtp_1
X_10456_ _10466_/CLK line[83] VGND VGND VPWR VPWR _10456_/Q sky130_fd_sc_hd__dfxtp_1
X_13175_ _13174_/Q _13202_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_10387_ _10386_/Q _10402_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09626__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ _12130_/CLK line[93] VGND VGND VPWR VPWR _12127_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[10\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12052__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12057_ _12057_/A _12082_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13726__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11008_ _11002_/CLK line[94] VGND VGND VPWR VPWR _11008_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06050__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11891__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06985__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].CGAND _13931_/X wr VGND VGND VPWR VPWR OVHB\[27\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA_OVHB\[27\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09361__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12959_ _12958_/Q _12992_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05500_ _05500_/CLK _05501_/X VGND VGND VPWR VPWR _05476_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10300__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06480_ _06480_/CLK _06481_/X VGND VGND VPWR VPWR _06464_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_53_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05431_ _13908_/X wr VGND VGND VPWR VPWR _05431_/X sky130_fd_sc_hd__and2_1
X_08150_ _08134_/CLK line[53] VGND VGND VPWR VPWR _08150_/Q sky130_fd_sc_hd__dfxtp_1
X_05362_ _13908_/X VGND VGND VPWR VPWR _05362_/Y sky130_fd_sc_hd__inv_2
X_07101_ _07101_/A _07112_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12227__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08081_ _08080_/Q _08092_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_05293_ _05299_/CLK line[32] VGND VGND VPWR VPWR _05293_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11131__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[9\].TOBUF OVHB\[18\].VALID\[9\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[4\].FF OVHB\[24\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[24\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09386__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07032_ _07030_/CLK line[54] VGND VGND VPWR VPWR _07032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06225__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09536__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08983_ _08982_/Q _09002_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13058__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07934_ _07946_/CLK line[82] VGND VGND VPWR VPWR _07934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07865_ _07865_/A _07882_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09604_ _09626_/CLK line[92] VGND VGND VPWR VPWR _09604_/Q sky130_fd_sc_hd__dfxtp_1
X_06816_ _06802_/CLK line[83] VGND VGND VPWR VPWR _06816_/Q sky130_fd_sc_hd__dfxtp_1
X_07796_ _07788_/CLK line[19] VGND VGND VPWR VPWR _07796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_MUX.MUX\[18\]_A0 _11435_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06747_ _06746_/Q _06762_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_09535_ _09534_/Q _09562_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[12\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11306__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09466_ _09482_/CLK line[29] VGND VGND VPWR VPWR _09466_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06678_ _06682_/CLK line[20] VGND VGND VPWR VPWR _06679_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05629_ _05628_/Q _05642_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_08417_ _08416_/Q _08442_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09397_ _09396_/Q _09422_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08348_ _08358_/CLK line[30] VGND VGND VPWR VPWR _08348_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08279_ _08279_/A _08302_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11041__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10310_ _10314_/CLK line[31] VGND VGND VPWR VPWR _10310_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06135__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11290_ _11302_/CLK line[95] VGND VGND VPWR VPWR _11290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10241_ _10240_/Q _10262_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10880__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05974__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08350__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10172_ _10188_/CLK line[81] VGND VGND VPWR VPWR _10173_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[6\].FF OVHB\[22\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[22\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[8\].TOBUF OVHB\[24\].VALID\[8\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[31\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13931_ _13934_/C _13934_/B _13933_/B _13934_/D VGND VGND VPWR VPWR _13931_/X sky130_fd_sc_hd__and4b_4
XFILLER_120_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[30\].VALID\[11\].FF OVHB\[30\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[30\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11066__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13862_ _13862_/A _13867_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12813_ _12803_/CLK line[9] VGND VGND VPWR VPWR _12814_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13793_ _13763_/CLK line[73] VGND VGND VPWR VPWR _13793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11216__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12744_ _12743_/Q _12747_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05214__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12675_/CLK _12676_/X VGND VGND VPWR VPWR _12667_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13431__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11626_ _11592_/A wr VGND VGND VPWR VPWR _11626_/X sky130_fd_sc_hd__and2_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _11592_/A VGND VGND VPWR VPWR _11557_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10508_ _10520_/CLK line[112] VGND VGND VPWR VPWR _10508_/Q sky130_fd_sc_hd__dfxtp_1
X_11488_ _11500_/CLK line[48] VGND VGND VPWR VPWR _11488_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10790__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13227_ _13213_/CLK line[70] VGND VGND VPWR VPWR _13227_/Q sky130_fd_sc_hd__dfxtp_1
X_10439_ _10438_/Q _10472_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[13\].FF OVHB\[20\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[20\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13158_ _13157_/Q _13167_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12109_ _12109_/CLK line[71] VGND VGND VPWR VPWR _12109_/Q sky130_fd_sc_hd__dfxtp_1
X_13089_ _13075_/CLK line[7] VGND VGND VPWR VPWR _13089_/Q sky130_fd_sc_hd__dfxtp_1
X_05980_ _05984_/CLK line[85] VGND VGND VPWR VPWR _05981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04931_ _04931_/A VGND VGND VPWR VPWR _04931_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[18\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13606__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07650_ _07644_/CLK line[95] VGND VGND VPWR VPWR _07650_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09091__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06601_ _06601_/A _06622_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07581_ _07581_/A _07602_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[11\].TOBUF OVHB\[3\].VALID\[11\].FF/Q OVHB\[3\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_09320_ _09320_/CLK line[90] VGND VGND VPWR VPWR _09320_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[8\].FF OVHB\[20\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[20\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06532_ _06528_/CLK line[81] VGND VGND VPWR VPWR _06532_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10030__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05124__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09251_ _09250_/Q _09282_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[7\].TOBUF OVHB\[30\].VALID\[7\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_06463_ _06462_/Q _06482_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10965__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08202_ _08208_/CLK line[91] VGND VGND VPWR VPWR _08202_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04963__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05414_ _05424_/CLK line[82] VGND VGND VPWR VPWR _05414_/Q sky130_fd_sc_hd__dfxtp_1
X_09182_ _09200_/CLK line[27] VGND VGND VPWR VPWR _09182_/Q sky130_fd_sc_hd__dfxtp_1
X_06394_ _06408_/CLK line[18] VGND VGND VPWR VPWR _06395_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[0\].TOBUF OVHB\[8\].VALID\[0\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08133_ _08132_/Q _08162_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
X_05345_ _05344_/Q _05362_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_08064_ _08070_/CLK line[28] VGND VGND VPWR VPWR _08064_/Q sky130_fd_sc_hd__dfxtp_1
X_05276_ _05278_/CLK line[19] VGND VGND VPWR VPWR _05276_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11796__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07015_ _07014_/Q _07042_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09266__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10205__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08966_ _13923_/X wr VGND VGND VPWR VPWR _08966_/X sky130_fd_sc_hd__and2_1
XOVHB\[17\].INV _13962_/X VGND VGND VPWR VPWR OVHB\[17\].INV/Y sky130_fd_sc_hd__inv_2
X_07917_ _13920_/X VGND VGND VPWR VPWR _07917_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08897_ _13923_/X VGND VGND VPWR VPWR _08897_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12420__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07848_ _07854_/CLK line[48] VGND VGND VPWR VPWR _07848_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07514__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[9\].FF OVHB\[19\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[19\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07779_ _07778_/Q _07812_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_09518_ _09518_/A _09527_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07811__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10790_ _10804_/CLK line[122] VGND VGND VPWR VPWR _10790_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _09427_/CLK line[7] VGND VGND VPWR VPWR _09450_/A sky130_fd_sc_hd__dfxtp_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12460_ _12459_/Q _12467_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[10\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11411_ _11395_/CLK line[8] VGND VGND VPWR VPWR _11411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12391_ _12387_/CLK line[72] VGND VGND VPWR VPWR _12391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11342_ _11341_/Q _11347_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11273_ _11251_/CLK line[73] VGND VGND VPWR VPWR _11273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10224_ _10223_/Q _10227_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_13012_ _13011_/Q _13027_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08080__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10155_ _10155_/CLK _10156_/X VGND VGND VPWR VPWR _10145_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09904__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10086_ _10192_/A wr VGND VGND VPWR VPWR _10086_/X sky130_fd_sc_hd__and2_1
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12330__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[3\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13914_ A[4] VGND VGND VPWR VPWR _13922_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13845_ _13845_/CLK line[111] VGND VGND VPWR VPWR _13846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[10\].CG clk OVHB\[10\].CGAND/X VGND VGND VPWR VPWR OVHB\[10\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_13776_ _13776_/A _13797_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_10988_ _10987_/Q _10997_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12727_ _12741_/CLK line[97] VGND VGND VPWR VPWR _12727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13161__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05879__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[13\].TOBUF OVHB\[26\].VALID\[13\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08255__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _12657_/Q _12677_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11609_ _11605_/CLK line[98] VGND VGND VPWR VPWR _11609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12589_ _12601_/CLK line[34] VGND VGND VPWR VPWR _12589_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05130_ _05122_/CLK line[95] VGND VGND VPWR VPWR _05130_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05061_ _05060_/Q _05082_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12505__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06503__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08820_ _08819_/Q _08827_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09814__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08751_ _08749_/CLK line[72] VGND VGND VPWR VPWR _08752_/A sky130_fd_sc_hd__dfxtp_1
X_05963_ _05962_/Q _05992_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[5\].TOBUF OVHB\[6\].VALID\[5\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13336__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07702_ _07702_/A _07707_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13914__A A[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05894_ _05902_/CLK line[60] VGND VGND VPWR VPWR _05894_/Q sky130_fd_sc_hd__dfxtp_1
X_08682_ _08682_/A _08687_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07633_ _07633_/CLK line[73] VGND VGND VPWR VPWR _07633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[23\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07564_ _07563_/Q _07567_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[15\]_A3 _13566_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06515_ _06515_/CLK _06516_/X VGND VGND VPWR VPWR _06489_/CLK sky130_fd_sc_hd__dlclkp_1
X_09303_ _09307_/CLK line[68] VGND VGND VPWR VPWR _09303_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05432__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10695__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07495_ _07495_/CLK _07496_/X VGND VGND VPWR VPWR _07467_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_16_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13071__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05789__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05151__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06446_ _06551_/A wr VGND VGND VPWR VPWR _06446_/X sky130_fd_sc_hd__and2_1
X_09234_ _09233_/Q _09247_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08165__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09165_ _09147_/CLK line[5] VGND VGND VPWR VPWR _09165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06377_ _06551_/A VGND VGND VPWR VPWR _06377_/Y sky130_fd_sc_hd__inv_2
X_08116_ _08115_/Q _08127_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_05328_ _05332_/CLK line[48] VGND VGND VPWR VPWR _05328_/Q sky130_fd_sc_hd__dfxtp_1
X_09096_ _09095_/Q _09107_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_08047_ _08033_/CLK line[6] VGND VGND VPWR VPWR _08047_/Q sky130_fd_sc_hd__dfxtp_1
X_05259_ _05258_/Q _05292_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06413__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13096__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05029__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09998_ _09997_/Q _10017_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05607__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08949_ _08947_/CLK line[34] VGND VGND VPWR VPWR _08949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13246__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05326__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11960_ _11959_/Q _11977_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07244__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10911_ _10903_/CLK line[35] VGND VGND VPWR VPWR _10911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11891_ _11901_/CLK line[99] VGND VGND VPWR VPWR _11891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13630_ _13629_/Q _13657_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_10842_ _10842_/A _10857_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13561_ _13559_/CLK line[109] VGND VGND VPWR VPWR _13561_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].CG clk OVHB\[5\].CGAND/X VGND VGND VPWR VPWR OVHB\[5\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_10773_ _10783_/CLK line[100] VGND VGND VPWR VPWR _10773_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[24\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[0\].TOBUF OVHB\[13\].VALID\[0\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_12512_ _12511_/Q _12537_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13492_ _13491_/Q _13517_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12443_ _12449_/CLK line[110] VGND VGND VPWR VPWR _12443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08803__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12374_ _12374_/A _12397_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11325_ _11343_/CLK line[111] VGND VGND VPWR VPWR _11326_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07419__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11256_ _11255_/Q _11277_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[19\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06901__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10207_ _10217_/CLK line[97] VGND VGND VPWR VPWR _10208_/A sky130_fd_sc_hd__dfxtp_1
X_11187_ _11191_/CLK line[33] VGND VGND VPWR VPWR _11188_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10138_ _10137_/Q _10157_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12060__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10069_ _10073_/CLK line[34] VGND VGND VPWR VPWR _10069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07154__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12995__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06993__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13828_ _13822_/CLK line[89] VGND VGND VPWR VPWR _13829_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13759_ _13758_/Q _13762_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06300_ _06299_/Q _06307_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
X_07280_ _07279_/Q _07287_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05402__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06231_ _06223_/CLK line[72] VGND VGND VPWR VPWR _06231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06162_ _06161_/Q _06167_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VOBUF OVHB\[15\].V/Q OVHB\[15\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XFILLER_102_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[13\].CGAND_A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[19\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _07915_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05113_ _05093_/CLK line[73] VGND VGND VPWR VPWR _05113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12235__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06093_ _06077_/CLK line[9] VGND VGND VPWR VPWR _06093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07329__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09921_ _09925_/CLK line[109] VGND VGND VPWR VPWR _09921_/Q sky130_fd_sc_hd__dfxtp_1
X_05044_ _05043_/Q _05047_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06233__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09852_ _09851_/Q _09877_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09544__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08803_ _08823_/CLK line[110] VGND VGND VPWR VPWR _08803_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04918__A2 _04918_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09783_ _09793_/CLK line[46] VGND VGND VPWR VPWR _09783_/Q sky130_fd_sc_hd__dfxtp_1
X_06995_ _07001_/CLK line[37] VGND VGND VPWR VPWR _06995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09841__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08734_ _08733_/Q _08757_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_05946_ _05946_/A _05957_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08665_ _08663_/CLK line[47] VGND VGND VPWR VPWR _08665_/Q sky130_fd_sc_hd__dfxtp_1
X_05877_ _05871_/CLK line[38] VGND VGND VPWR VPWR _05877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07616_ _07616_/A _07637_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
X_08596_ _08595_/Q _08617_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07547_ _07539_/CLK line[33] VGND VGND VPWR VPWR _07548_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07478_ _07477_/Q _07497_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06408__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09217_ _09241_/CLK line[43] VGND VGND VPWR VPWR _09217_/Q sky130_fd_sc_hd__dfxtp_1
X_06429_ _06421_/CLK line[34] VGND VGND VPWR VPWR _06429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09719__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09148_ _09147_/Q _09177_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09079_ _09085_/CLK line[108] VGND VGND VPWR VPWR _09080_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _11109_/Q _11137_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06143__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12090_ _12089_/Q _12117_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11984__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[6\].FF OVHB\[8\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[8\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11041_ _11063_/CLK line[109] VGND VGND VPWR VPWR _11041_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[18\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _07530_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_104_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05982__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[11\].VALID\[5\].TOBUF OVHB\[11\].VALID\[5\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_76_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12992_ _12992_/A VGND VGND VPWR VPWR _12992_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11943_ _11945_/CLK line[0] VGND VGND VPWR VPWR _11943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11874_ _11873_/Q _11907_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_13613_ _13612_/Q _13622_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_10825_ _10843_/CLK line[10] VGND VGND VPWR VPWR _10825_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11224__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11802__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13544_ _13528_/CLK line[87] VGND VGND VPWR VPWR _13544_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06318__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10756_ _10755_/Q _10787_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[25\].VALID\[13\].FF OVHB\[25\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[25\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11521__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13475_ _13475_/A _13482_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10687_ _10707_/CLK line[75] VGND VGND VPWR VPWR _10687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08533__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[5\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12426_ _12414_/CLK line[88] VGND VGND VPWR VPWR _12427_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[22\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12357_ _12357_/A _12362_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
X_11308_ _11302_/CLK line[89] VGND VGND VPWR VPWR _11309_/A sky130_fd_sc_hd__dfxtp_1
X_12288_ _12268_/CLK line[25] VGND VGND VPWR VPWR _12288_/Q sky130_fd_sc_hd__dfxtp_1
X_11239_ _11238_/Q _11242_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05892__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05800_ _05800_/A _05817_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_06780_ _06779_/Q _06797_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05731_ _05739_/CLK line[99] VGND VGND VPWR VPWR _05731_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07462__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[8\].FF OVHB\[6\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[6\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13614__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08450_ _08449_/Q _08477_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_05662_ _05661_/Q _05677_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07181__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08708__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07401_ _07393_/CLK line[109] VGND VGND VPWR VPWR _07401_/Q sky130_fd_sc_hd__dfxtp_1
X_08381_ _08383_/CLK line[45] VGND VGND VPWR VPWR _08381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[16\].VALID\[11\].TOBUF OVHB\[16\].VALID\[11\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05593_ _05575_/CLK line[36] VGND VGND VPWR VPWR _05593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07332_ _07331_/Q _07357_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05132__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07263_ _07267_/CLK line[46] VGND VGND VPWR VPWR _07263_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10973__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09002_ _13923_/X VGND VGND VPWR VPWR _09002_/Y sky130_fd_sc_hd__inv_2
X_06214_ _06213_/Q _06237_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08443__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04971__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07194_ _07193_/Q _07217_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06145_ _06147_/CLK line[47] VGND VGND VPWR VPWR _06146_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07059__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07637__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06076_ _06075_/Q _06097_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_05027_ _05041_/CLK line[33] VGND VGND VPWR VPWR _05027_/Q sky130_fd_sc_hd__dfxtp_1
X_09904_ _09908_/CLK line[87] VGND VGND VPWR VPWR _09904_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07356__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06898__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09274__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09835_ _09834_/Q _09842_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10213__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09766_ _09760_/CLK line[24] VGND VGND VPWR VPWR _09766_/Q sky130_fd_sc_hd__dfxtp_1
X_06978_ _06978_/A _07007_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05307__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08717_ _08717_/A _08722_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05929_ _05929_/CLK line[76] VGND VGND VPWR VPWR _05929_/Q sky130_fd_sc_hd__dfxtp_1
X_09697_ _09696_/Q _09702_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13524__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08618__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08648_ _08646_/CLK line[25] VGND VGND VPWR VPWR _08648_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07522__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _08579_/A _08582_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[22\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _10610_/CLK _10611_/X VGND VGND VPWR VPWR _10594_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _11590_/CLK _11591_/X VGND VGND VPWR VPWR _11588_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _13931_/X wr VGND VGND VPWR VPWR _10541_/X sky130_fd_sc_hd__and2_1
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _13254_/CLK line[85] VGND VGND VPWR VPWR _13260_/Q sky130_fd_sc_hd__dfxtp_1
X_10472_ _13931_/X VGND VGND VPWR VPWR _10472_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08931__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ _12210_/Q _12222_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[28\]_A2 _06525_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13191_ _13190_/Q _13202_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12142_ _12130_/CLK line[86] VGND VGND VPWR VPWR _12142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12603__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ _12073_/A _12082_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09184__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11024_ _11002_/CLK line[87] VGND VGND VPWR VPWR _11025_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10123__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12975_ _12974_/Q _12992_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_11926_ _11934_/CLK line[115] VGND VGND VPWR VPWR _11927_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07432__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[0\].FF OVHB\[15\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[15\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11857_ _11856_/Q _11872_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[3\] _11402_/Z _05592_/Z _13502_/Z _13572_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[3] sky130_fd_sc_hd__mux4_1
XANTENNA__06048__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10808_ _10804_/CLK line[116] VGND VGND VPWR VPWR _10808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11788_ _11776_/CLK line[52] VGND VGND VPWR VPWR _11788_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11889__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09002__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13527_ _13526_/Q _13552_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_10739_ _10739_/A _10752_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09359__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08263__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13458_ _13468_/CLK line[62] VGND VGND VPWR VPWR _13458_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].CGAND _09352_/A wr VGND VGND VPWR VPWR OVHB\[23\].CGAND/X sky130_fd_sc_hd__and2_4
X_12409_ _12408_/Q _12432_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13389_ _13388_/Q _13412_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12513__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07950_ _07950_/CLK _07951_/X VGND VGND VPWR VPWR _07946_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07607__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06511__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06901_ _06832_/A wr VGND VGND VPWR VPWR _06901_/X sky130_fd_sc_hd__and2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[20\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07881_ _13920_/X wr VGND VGND VPWR VPWR _07881_/X sky130_fd_sc_hd__and2_1
XANTENNA__11129__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09620_ _09626_/CLK line[85] VGND VGND VPWR VPWR _09621_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06832_ _06832_/A VGND VGND VPWR VPWR _06832_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10611__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09822__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09551_ _09550_/Q _09562_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[5\].TOBUF OVHB\[18\].VALID\[5\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06763_ _06775_/CLK line[64] VGND VGND VPWR VPWR _06763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[21\].VALID\[11\].FF OVHB\[21\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[21\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08502_ _08480_/CLK line[86] VGND VGND VPWR VPWR _08503_/A sky130_fd_sc_hd__dfxtp_1
X_05714_ _05713_/Q _05747_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08438__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06694_ _06693_/Q _06727_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_09482_ _09482_/CLK line[22] VGND VGND VPWR VPWR _09482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08433_ _08433_/A _08442_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_05645_ _05671_/CLK line[74] VGND VGND VPWR VPWR _05645_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05576_ _05575_/Q _05607_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08364_ _08358_/CLK line[23] VGND VGND VPWR VPWR _08364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07315_ _07314_/Q _07322_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_08295_ _08294_/Q _08302_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05797__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08173__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07246_ _07232_/CLK line[24] VGND VGND VPWR VPWR _07246_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[2\].FF OVHB\[13\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[13\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07177_ _07176_/Q _07182_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[6\].FF OVHB\[30\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[30\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06128_ _06108_/CLK line[25] VGND VGND VPWR VPWR _06128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06271__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06059_ _06059_/A _06062_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[11\].VALID\[13\].FF OVHB\[11\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[11\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06421__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[27\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11039__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09818_ _09834_/CLK line[62] VGND VGND VPWR VPWR _09819_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05037__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10878__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09749_ _09748_/Q _09772_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13254__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13832__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12760_ _12774_/CLK line[127] VGND VGND VPWR VPWR _12760_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11710_/Q _11732_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13551__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12690_/Q _12712_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11636_/CLK line[113] VGND VGND VPWR VPWR _11643_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06446__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[4\].TOBUF OVHB\[24\].VALID\[4\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _11573_/A _11592_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11502__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13308_/CLK line[123] VGND VGND VPWR VPWR _13313_/A sky130_fd_sc_hd__dfxtp_1
X_10524_ _10520_/CLK line[114] VGND VGND VPWR VPWR _10524_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VALID\[7\].FF OVHB\[29\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[29\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10118__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13243_ _13242_/Q _13272_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_10455_ _10454_/Q _10472_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08811__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13174_ _13194_/CLK line[60] VGND VGND VPWR VPWR _13174_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _13830_/CLK sky130_fd_sc_hd__clkbuf_4
X_10386_ _10384_/CLK line[51] VGND VGND VPWR VPWR _10386_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13429__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12125_ _12124_/Q _12152_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[19\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[4\].FF OVHB\[11\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[11\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09492__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13726__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12056_ _12072_/CLK line[61] VGND VGND VPWR VPWR _12057_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11007_ _11006_/Q _11032_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10788__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12958_ _12962_/CLK line[80] VGND VGND VPWR VPWR _12958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07162__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11909_ _11908_/Q _11942_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12889_ _12888_/Q _12922_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05430_ _05430_/CLK _05431_/X VGND VGND VPWR VPWR _05424_/CLK sky130_fd_sc_hd__dlclkp_1
X_05361_ _13908_/X wr VGND VGND VPWR VPWR _05361_/X sky130_fd_sc_hd__and2_1
XANTENNA__09089__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07100_ _07098_/CLK line[85] VGND VGND VPWR VPWR _07101_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09667__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08080_ _08070_/CLK line[21] VGND VGND VPWR VPWR _08080_/Q sky130_fd_sc_hd__dfxtp_1
X_05292_ _13908_/X VGND VGND VPWR VPWR _05292_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05410__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07031_ _07031_/A _07042_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10028__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09386__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12243__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08982_ _08972_/CLK line[49] VGND VGND VPWR VPWR _08982_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07337__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[3\].TOBUF OVHB\[30\].VALID\[3\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_114_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[27\].VALID\[9\].FF OVHB\[27\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[27\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07933_ _07932_/Q _07952_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[8\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _13445_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_29_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07864_ _07854_/CLK line[50] VGND VGND VPWR VPWR _07865_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09552__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09603_ _09602_/Q _09632_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_06815_ _06814_/Q _06832_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_07795_ _07794_/Q _07812_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09534_ _09554_/CLK line[60] VGND VGND VPWR VPWR _09534_/Q sky130_fd_sc_hd__dfxtp_1
X_06746_ _06740_/CLK line[51] VGND VGND VPWR VPWR _06746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[18\]_A1 _13465_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09465_ _09464_/Q _09492_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06677_ _06677_/A _06692_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13802__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08416_ _08410_/CLK line[61] VGND VGND VPWR VPWR _08416_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05628_ _05632_/CLK line[52] VGND VGND VPWR VPWR _05628_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09396_ _09414_/CLK line[125] VGND VGND VPWR VPWR _09396_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07800__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08347_ _08346_/Q _08372_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12418__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05559_ _05558_/Q _05572_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ _08282_/CLK line[126] VGND VGND VPWR VPWR _08279_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07229_ _07228_/Q _07252_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09727__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[28\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _10785_/CLK sky130_fd_sc_hd__clkbuf_4
X_10240_ _10248_/CLK line[127] VGND VGND VPWR VPWR _10240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12153__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10171_ _10171_/A _10192_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06151__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11992__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11347__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ _13934_/C _13933_/B _13934_/B _13934_/D VGND VGND VPWR VPWR _10192_/A sky130_fd_sc_hd__and4bb_4
XFILLER_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[9\].TOBUF OVHB\[22\].VALID\[9\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09462__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13861_ _13845_/CLK line[104] VGND VGND VPWR VPWR _13862_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11066__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12812_ _12812_/A _12817_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08078__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ _13792_/A _13797_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[13\].TOBUF OVHB\[6\].VALID\[13\].FF/Q OVHB\[6\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_12743_ _12741_/CLK line[105] VGND VGND VPWR VPWR _12743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12673_/Q _12677_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11625_ _11625_/CLK _11626_/X VGND VGND VPWR VPWR _11605_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11232__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06326__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _11592_/A wr VGND VGND VPWR VPWR _11556_/X sky130_fd_sc_hd__and2_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ _13931_/X VGND VGND VPWR VPWR _10507_/Y sky130_fd_sc_hd__inv_2
X_11487_ _11592_/A VGND VGND VPWR VPWR _11487_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09637__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08541__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13226_ _13225_/Q _13237_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_10438_ _10466_/CLK line[80] VGND VGND VPWR VPWR _10438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13159__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ _13163_/CLK line[38] VGND VGND VPWR VPWR _13157_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12641__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10369_ _10368_/Q _10402_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_12108_ _12107_/Q _12117_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
X_13088_ _13088_/A _13097_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[27\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _10400_/CLK sky130_fd_sc_hd__clkbuf_4
X_04930_ _04923_/X _04926_/Y _04928_/X _04929_/X VGND VGND VPWR VPWR _04931_/A sky130_fd_sc_hd__or4_4
X_12039_ _12019_/CLK line[39] VGND VGND VPWR VPWR _12039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[31\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11407__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06600_ _06596_/CLK line[127] VGND VGND VPWR VPWR _06601_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07580_ _07572_/CLK line[63] VGND VGND VPWR VPWR _07581_/A sky130_fd_sc_hd__dfxtp_1
X_06531_ _06530_/Q _06552_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09250_ _09256_/CLK line[58] VGND VGND VPWR VPWR _09250_/Q sky130_fd_sc_hd__dfxtp_1
X_06462_ _06464_/CLK line[49] VGND VGND VPWR VPWR _06462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08716__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08201_ _08200_/Q _08232_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_05413_ _05413_/A _05432_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_06393_ _06393_/A _06412_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
X_09181_ _09180_/Q _09212_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11142__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12816__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08132_ _08134_/CLK line[59] VGND VGND VPWR VPWR _08132_/Q sky130_fd_sc_hd__dfxtp_1
X_05344_ _05332_/CLK line[50] VGND VGND VPWR VPWR _05344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[6\].VALID\[1\].TOBUF OVHB\[6\].VALID\[1\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05140__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10981__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05275_ _05275_/A _05292_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
X_08063_ _08063_/A _08092_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07014_ _07030_/CLK line[60] VGND VGND VPWR VPWR _07014_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08451__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13069__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07067__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08965_ _08965_/CLK _08966_/X VGND VGND VPWR VPWR _08947_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[12\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07916_ _13920_/X wr VGND VGND VPWR VPWR _07916_/X sky130_fd_sc_hd__and2_1
XFILLER_116_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08896_ _13923_/X wr VGND VGND VPWR VPWR _08896_/X sky130_fd_sc_hd__and2_1
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07847_ _13920_/X VGND VGND VPWR VPWR _07847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11317__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10221__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[26\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _10015_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08476__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07778_ _07788_/CLK line[16] VGND VGND VPWR VPWR _07778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05315__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09517_ _09507_/CLK line[38] VGND VGND VPWR VPWR _09518_/A sky130_fd_sc_hd__dfxtp_1
X_06729_ _06728_/Q _06762_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13532__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[16\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _07145_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _09447_/Q _09457_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08626__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XMUX.MUX\[21\] _10881_/Z _10391_/Z _13541_/Z _07171_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[21] sky130_fd_sc_hd__mux4_1
XANTENNA__12148__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09379_ _09365_/CLK line[103] VGND VGND VPWR VPWR _09379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11410_ _11409_/Q _11417_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05050__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12390_ _12389_/Q _12397_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11341_ _11343_/CLK line[104] VGND VGND VPWR VPWR _11341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[2\].VALID\[13\].FF OVHB\[2\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[2\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11272_ _11271_/Q _11277_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[27\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13011_ _12999_/CLK line[99] VGND VGND VPWR VPWR _13011_/Q sky130_fd_sc_hd__dfxtp_1
X_10223_ _10217_/CLK line[105] VGND VGND VPWR VPWR _10223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04939__B1 A_h[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10154_ _10154_/A _10157_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13707__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10085_ _10085_/CLK _10086_/X VGND VGND VPWR VPWR _10073_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09192__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ _13909_/C _13909_/B _13905_/X _13909_/D VGND VGND VPWR VPWR _06832_/A sky130_fd_sc_hd__and4_4
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[22\].VALID\[14\].TOBUF OVHB\[22\].VALID\[14\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__10131__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13844_ _13843_/Q _13867_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05225__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13775_ _13763_/CLK line[79] VGND VGND VPWR VPWR _13776_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10987_ _10977_/CLK line[70] VGND VGND VPWR VPWR _10987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ _12725_/Q _12747_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07440__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12058__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ _12667_/CLK line[65] VGND VGND VPWR VPWR _12657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11608_/A _11627_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06056__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[15\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _06760_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[14\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[1\].FF OVHB\[0\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[0\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12588_ _12588_/A _12607_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11897__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11539_ _11535_/CLK line[66] VGND VGND VPWR VPWR _11540_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10156__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09367__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05060_ _05058_/CLK line[63] VGND VGND VPWR VPWR _05060_/Q sky130_fd_sc_hd__dfxtp_1
X_13209_ _13213_/CLK line[76] VGND VGND VPWR VPWR _13209_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10306__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[11\].FF OVHB\[26\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[26\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12521__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08750_ _08749_/Q _08757_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05962_ _05984_/CLK line[91] VGND VGND VPWR VPWR _05962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07615__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07701_ _07679_/CLK line[104] VGND VGND VPWR VPWR _07702_/A sky130_fd_sc_hd__dfxtp_1
X_08681_ _08663_/CLK line[40] VGND VGND VPWR VPWR _08682_/A sky130_fd_sc_hd__dfxtp_1
X_05893_ _05893_/A _05922_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[4\].VALID\[6\].TOBUF OVHB\[4\].VALID\[6\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VOBUF OVHB\[11\].V/Q OVHB\[11\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_07632_ _07631_/Q _07637_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[9\].TOBUF OVHB\[29\].VALID\[9\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09830__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07563_ _07539_/CLK line[41] VGND VGND VPWR VPWR _07563_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[23\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09302_ _09301_/Q _09317_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06514_ _06513_/Q _06517_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07494_ _07493_/Q _07497_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09233_ _09241_/CLK line[36] VGND VGND VPWR VPWR _09233_/Q sky130_fd_sc_hd__dfxtp_1
X_06445_ _06445_/CLK _06446_/X VGND VGND VPWR VPWR _06421_/CLK sky130_fd_sc_hd__dlclkp_1
X_09164_ _09163_/Q _09177_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_06376_ _06551_/A wr VGND VGND VPWR VPWR _06376_/X sky130_fd_sc_hd__and2_1
XFILLER_119_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[16\].VALID\[13\].FF OVHB\[16\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[16\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08115_ _08113_/CLK line[37] VGND VGND VPWR VPWR _08115_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[11\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05327_ _13908_/X VGND VGND VPWR VPWR _05327_/Y sky130_fd_sc_hd__inv_2
X_09095_ _09085_/CLK line[101] VGND VGND VPWR VPWR _09095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08181__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08046_ _08045_/Q _08057_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_05258_ _05278_/CLK line[16] VGND VGND VPWR VPWR _05258_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[14\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _06375_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13377__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05189_ _05188_/Q _05222_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13096__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ _10011_/CLK line[1] VGND VGND VPWR VPWR _09997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08948_ _08947_/Q _08967_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08879_ _08869_/CLK line[2] VGND VGND VPWR VPWR _08879_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11047__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10910_ _10909_/Q _10927_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11890_ _11890_/A _11907_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[4\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09740__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10841_ _10843_/CLK line[3] VGND VGND VPWR VPWR _10842_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10886__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13262__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13560_ _13560_/A _13587_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08356__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10772_ _10771_/Q _10787_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[30\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12511_ _12523_/CLK line[13] VGND VGND VPWR VPWR _12511_/Q sky130_fd_sc_hd__dfxtp_1
X_13491_ _13497_/CLK line[77] VGND VGND VPWR VPWR _13491_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[1\].TOBUF OVHB\[11\].VALID\[1\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_12442_ _12441_/Q _12467_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12373_ _12387_/CLK line[78] VGND VGND VPWR VPWR _12374_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11510__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11324_ _11323_/Q _11347_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06604__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11255_ _11251_/CLK line[79] VGND VGND VPWR VPWR _11255_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06901__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09915__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10206_ _10205_/Q _10227_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_11186_ _11185_/Q _11207_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13437__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10137_ _10145_/CLK line[65] VGND VGND VPWR VPWR _10137_/Q sky130_fd_sc_hd__dfxtp_1
X_10068_ _10068_/A _10087_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10796__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13827_ _13827_/A _13832_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13172__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13758_ _13746_/CLK line[57] VGND VGND VPWR VPWR _13758_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07170__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12709_ _12708_/Q _12712_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13689_ _13688_/Q _13692_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06230_ _06230_/A _06237_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[16\].INV _13961_/Y VGND VGND VPWR VPWR OVHB\[16\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[29\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06161_ _06147_/CLK line[40] VGND VGND VPWR VPWR _06161_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09097__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11420__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05112_ _05112_/A _05117_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_06092_ _06091_/Q _06097_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_09920_ _09919_/Q _09947_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
X_05043_ _05041_/CLK line[41] VGND VGND VPWR VPWR _05043_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10036__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].CGAND_A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09851_ _09849_/CLK line[77] VGND VGND VPWR VPWR _09851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13347__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08802_ _08801_/Q _08827_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12251__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04969__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13925__A A[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09782_ _09782_/A _09807_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_06994_ _06994_/A _07007_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07345__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08733_ _08749_/CLK line[78] VGND VGND VPWR VPWR _08733_/Q sky130_fd_sc_hd__dfxtp_1
X_05945_ _05929_/CLK line[69] VGND VGND VPWR VPWR _05946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08664_ _08664_/A _08687_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_05876_ _05875_/Q _05887_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].CGAND _07672_/A wr VGND VGND VPWR VPWR OVHB\[18\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07615_ _07633_/CLK line[79] VGND VGND VPWR VPWR _07616_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08595_ _08609_/CLK line[15] VGND VGND VPWR VPWR _08595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[29\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _07545_/Q _07567_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07080__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ _07467_/CLK line[1] VGND VGND VPWR VPWR _07477_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13810__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09216_ _09215_/Q _09247_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
X_06428_ _06428_/A _06447_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08904__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09147_ _09147_/CLK line[11] VGND VGND VPWR VPWR _09147_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12426__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06359_ _06353_/CLK line[2] VGND VGND VPWR VPWR _06359_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09078_ _09077_/Q _09107_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_08029_ _08033_/CLK line[12] VGND VGND VPWR VPWR _08030_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11040_ _11040_/A _11067_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12161__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[23\].VALID\[0\].FF OVHB\[23\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[23\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07255__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12991_ _12992_/A wr VGND VGND VPWR VPWR _12991_/X sky130_fd_sc_hd__and2_1
X_11942_ _11872_/A VGND VGND VPWR VPWR _11942_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09470__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11873_ _11901_/CLK line[96] VGND VGND VPWR VPWR _11873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13612_ _13598_/CLK line[118] VGND VGND VPWR VPWR _13612_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[11\].FF OVHB\[12\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[12\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10824_ _10824_/A _10857_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08086__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05503__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[13\].TOBUF OVHB\[19\].VALID\[13\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_13543_ _13542_/Q _13552_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10755_ _10783_/CLK line[106] VGND VGND VPWR VPWR _10755_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12186__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[2\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13474_ _13468_/CLK line[55] VGND VGND VPWR VPWR _13475_/A sky130_fd_sc_hd__dfxtp_1
X_10686_ _10685_/Q _10717_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_12425_ _12425_/A _12432_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12336__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[5\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06334__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12356_ _12352_/CLK line[56] VGND VGND VPWR VPWR _12357_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[23\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _11306_/Q _11312_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_MUX.MUX\[13\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12287_ _12287_/A _12292_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09645__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11238_ _11216_/CLK line[57] VGND VGND VPWR VPWR _11238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11169_ _11168_/Q _11172_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[16\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[12\].TOBUF OVHB\[12\].VALID\[12\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_05730_ _05729_/Q _05747_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05661_ _05671_/CLK line[67] VGND VGND VPWR VPWR _05661_/Q sky130_fd_sc_hd__dfxtp_1
X_07400_ _07399_/Q _07427_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[2\].FF OVHB\[21\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[21\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08380_ _08380_/A _08407_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06509__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05592_ _05591_/Q _05607_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_07331_ _07327_/CLK line[77] VGND VGND VPWR VPWR _07331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[6\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _13060_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_32_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ _07261_/Q _07287_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_09001_ _13923_/X wr VGND VGND VPWR VPWR _09001_/X sky130_fd_sc_hd__and2_1
X_06213_ _06223_/CLK line[78] VGND VGND VPWR VPWR _06213_/Q sky130_fd_sc_hd__dfxtp_1
X_07193_ _07183_/CLK line[14] VGND VGND VPWR VPWR _07193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11150__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[1\].TOBUF OVHB\[18\].VALID\[1\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].CG clk OVHB\[23\].CGAND/X VGND VGND VPWR VPWR OVHB\[23\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_06144_ _06143_/Q _06167_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06244__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06075_ _06077_/CLK line[15] VGND VGND VPWR VPWR _06075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05026_ _05025_/Q _05047_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_09903_ _09902_/Q _09912_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13077__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09834_ _09834_/CLK line[55] VGND VGND VPWR VPWR _09834_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09765_ _09764_/Q _09772_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_06977_ _07001_/CLK line[43] VGND VGND VPWR VPWR _06978_/A sky130_fd_sc_hd__dfxtp_1
X_08716_ _08710_/CLK line[56] VGND VGND VPWR VPWR _08717_/A sky130_fd_sc_hd__dfxtp_1
X_05928_ _05927_/Q _05957_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_09696_ _09694_/CLK line[120] VGND VGND VPWR VPWR _09696_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08647_ _08646_/Q _08652_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_05859_ _05871_/CLK line[44] VGND VGND VPWR VPWR _05860_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11325__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06419__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ _08560_/CLK line[121] VGND VGND VPWR VPWR _08579_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05323__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ _07529_/A _07532_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13540__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[7\].VALID\[13\].FF OVHB\[7\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[7\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10540_ _10540_/CLK _10541_/X VGND VGND VPWR VPWR _10520_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08634__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[27\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ _13931_/X wr VGND VGND VPWR VPWR _10471_/X sky130_fd_sc_hd__and2_1
XANTENNA__08931__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[5\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _12675_/CLK sky130_fd_sc_hd__clkbuf_4
X_12210_ _12204_/CLK line[117] VGND VGND VPWR VPWR _12210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13190_ _13194_/CLK line[53] VGND VGND VPWR VPWR _13190_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[28\]_A3 _13595_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12141_ _12140_/Q _12152_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05993__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12072_ _12072_/CLK line[54] VGND VGND VPWR VPWR _12073_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11023_ _11023_/A _11032_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[24\].VALID\[0\].TOBUF OVHB\[24\].VALID\[0\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13715__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08809__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12974_ _12962_/CLK line[82] VGND VGND VPWR VPWR _12974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11925_ _11924_/Q _11942_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11856_ _11846_/CLK line[83] VGND VGND VPWR VPWR _11856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05233__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10807_ _10807_/A _10822_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_11787_ _11786_/Q _11802_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13450__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13526_ _13528_/CLK line[93] VGND VGND VPWR VPWR _13526_/Q sky130_fd_sc_hd__dfxtp_1
X_10738_ _10728_/CLK line[84] VGND VGND VPWR VPWR _10739_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[18\].VALID\[5\].FF OVHB\[18\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[18\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12066__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13457_ _13456_/Q _13482_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_10669_ _10668_/Q _10682_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_12408_ _12414_/CLK line[94] VGND VGND VPWR VPWR _12408_/Q sky130_fd_sc_hd__dfxtp_1
X_13388_ _13394_/CLK line[30] VGND VGND VPWR VPWR _13388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[0\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12339_ _12339_/A _12362_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06999__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].V OVHB\[1\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[1\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09375__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[4\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _12290_/CLK sky130_fd_sc_hd__clkbuf_4
X_06900_ _06900_/CLK _06901_/X VGND VGND VPWR VPWR _06892_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10314__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07880_ _07880_/CLK _07881_/X VGND VGND VPWR VPWR _07854_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05408__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06831_ _06832_/A wr VGND VGND VPWR VPWR _06831_/X sky130_fd_sc_hd__and2_1
XFILLER_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13625__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10611__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09550_ _09554_/CLK line[53] VGND VGND VPWR VPWR _09550_/Q sky130_fd_sc_hd__dfxtp_1
X_06762_ _06832_/A VGND VGND VPWR VPWR _06762_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07623__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[6\].TOBUF OVHB\[16\].VALID\[6\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_08501_ _08500_/Q _08512_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05713_ _05739_/CLK line[96] VGND VGND VPWR VPWR _05713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09481_ _09480_/Q _09492_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_06693_ _06711_/CLK line[32] VGND VGND VPWR VPWR _06693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08432_ _08410_/CLK line[54] VGND VGND VPWR VPWR _08433_/A sky130_fd_sc_hd__dfxtp_1
X_05644_ _05643_/Q _05677_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08363_ _08362_/Q _08372_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_05575_ _05575_/CLK line[42] VGND VGND VPWR VPWR _05575_/Q sky130_fd_sc_hd__dfxtp_1
X_07314_ _07292_/CLK line[55] VGND VGND VPWR VPWR _07314_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04982__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08294_ _08282_/CLK line[119] VGND VGND VPWR VPWR _08294_/Q sky130_fd_sc_hd__dfxtp_1
X_07245_ _07244_/Q _07252_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[24\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _09630_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_30_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07176_ _07170_/CLK line[120] VGND VGND VPWR VPWR _07176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06552__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06127_ _06126_/Q _06132_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12704__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04920__A2_N _04920_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06271__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09285__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[7\].FF OVHB\[16\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[16\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06058_ _06050_/CLK line[121] VGND VGND VPWR VPWR _06059_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05009_ _05008_/Q _05012_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04935__A2_N _04935_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09817_ _09817_/A _09842_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _09760_/CLK line[30] VGND VGND VPWR VPWR _09748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07533__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09679_ _09678_/Q _09702_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11055__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11706_/CLK line[31] VGND VGND VPWR VPWR _11710_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06149__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12708_/CLK line[95] VGND VGND VPWR VPWR _12690_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11641_ _11641_/A _11662_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06446__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05988__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[28\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _11588_/CLK line[81] VGND VGND VPWR VPWR _11573_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13310_/Q _13342_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10523_ _10522_/Q _10542_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[22\].VALID\[5\].TOBUF OVHB\[22\].VALID\[5\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13242_ _13254_/CLK line[91] VGND VGND VPWR VPWR _13242_/Q sky130_fd_sc_hd__dfxtp_1
X_10454_ _10466_/CLK line[82] VGND VGND VPWR VPWR _10454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13173_ _13172_/Q _13202_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12614__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10385_ _10384_/Q _10402_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07708__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12124_ _12130_/CLK line[92] VGND VGND VPWR VPWR _12124_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _09245_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06612__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[12\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12055_ _12054_/Q _12082_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09923__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11006_ _11002_/CLK line[93] VGND VGND VPWR VPWR _11006_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08539__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[9\].FF OVHB\[14\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[14\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[11\].FF OVHB\[3\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[3\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12957_ _12992_/A VGND VGND VPWR VPWR _12957_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11908_ _11934_/CLK line[112] VGND VGND VPWR VPWR _11908_/Q sky130_fd_sc_hd__dfxtp_1
X_12888_ _12902_/CLK line[48] VGND VGND VPWR VPWR _12888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11839_ _11839_/A _11872_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13180__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05898__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05360_ _05360_/CLK _05361_/X VGND VGND VPWR VPWR _05332_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08274__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13509_ _13497_/CLK line[71] VGND VGND VPWR VPWR _13509_/Q sky130_fd_sc_hd__dfxtp_1
X_05291_ _13908_/X wr VGND VGND VPWR VPWR _05291_/X sky130_fd_sc_hd__and2_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07030_ _07030_/CLK line[53] VGND VGND VPWR VPWR _07031_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06522__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08981_ _08980_/Q _09002_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10044__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07932_ _07946_/CLK line[81] VGND VGND VPWR VPWR _07932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05138__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07863_ _07863_/A _07882_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10979__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13355__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09602_ _09626_/CLK line[91] VGND VGND VPWR VPWR _09602_/Q sky130_fd_sc_hd__dfxtp_1
X_06814_ _06802_/CLK line[82] VGND VGND VPWR VPWR _06814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08449__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07794_ _07788_/CLK line[18] VGND VGND VPWR VPWR _07794_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07353__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09533_ _09532_/Q _09562_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06745_ _06744_/Q _06762_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[12\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _05990_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_MUX.MUX\[18\]_A2 _07095_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09464_ _09482_/CLK line[28] VGND VGND VPWR VPWR _09464_/Q sky130_fd_sc_hd__dfxtp_1
X_06676_ _06682_/CLK line[19] VGND VGND VPWR VPWR _06677_/A sky130_fd_sc_hd__dfxtp_1
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _08414_/Q _08442_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_05627_ _05626_/Q _05642_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_09395_ _09394_/Q _09422_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11603__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08346_ _08358_/CLK line[29] VGND VGND VPWR VPWR _08346_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05558_ _05568_/CLK line[20] VGND VGND VPWR VPWR _05558_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05601__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10219__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08277_ _08276_/Q _08302_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_05489_ _05488_/Q _05502_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07228_ _07232_/CLK line[30] VGND VGND VPWR VPWR _07228_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08912__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07159_ _07158_/Q _07182_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[25\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07528__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10170_ _10188_/CLK line[95] VGND VGND VPWR VPWR _10171_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[0\].FF OVHB\[9\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[9\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[11\].TOBUF OVHB\[29\].VALID\[11\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05048__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[14\].TOBUF OVHB\[2\].VALID\[14\].FF/Q OVHB\[2\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_86_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[17\].VALID\[11\].FF OVHB\[17\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[17\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13860_ _13860_/A _13867_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07263__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12811_ _12803_/CLK line[8] VGND VGND VPWR VPWR _12812_/A sky130_fd_sc_hd__dfxtp_1
X_13791_ _13763_/CLK line[72] VGND VGND VPWR VPWR _13792_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12742_ _12741_/Q _12747_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05361__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12667_/CLK line[73] VGND VGND VPWR VPWR _12673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _05605_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_MUX.MUX\[0\]_A0 _06904_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11623_/Q _11627_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05511__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10129__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11555_ _11555_/CLK _11556_/X VGND VGND VPWR VPWR _11535_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10506_ _13931_/X wr VGND VGND VPWR VPWR _10506_/X sky130_fd_sc_hd__and2_1
X_11486_ _11592_/A wr VGND VGND VPWR VPWR _11486_/X sky130_fd_sc_hd__and2_1
XOVHB\[22\].VALID\[10\].TOBUF OVHB\[22\].VALID\[10\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_87_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13225_ _13213_/CLK line[69] VGND VGND VPWR VPWR _13225_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12344__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10437_ _13931_/X VGND VGND VPWR VPWR _10437_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12922__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07438__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13156_ _13155_/Q _13167_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
X_10368_ _10384_/CLK line[48] VGND VGND VPWR VPWR _10368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12641__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _12109_/CLK line[70] VGND VGND VPWR VPWR _12107_/Q sky130_fd_sc_hd__dfxtp_1
X_13087_ _13075_/CLK line[6] VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__dfxtp_1
X_10299_ _10298_/Q _10332_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09653__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05536__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12038_ _12037_/Q _12047_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[6\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[2\].FF OVHB\[7\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[7\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13989_ _13990_/A _13990_/B _13982_/X _13990_/D VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__and4b_4
X_06530_ _06528_/CLK line[95] VGND VGND VPWR VPWR _06530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07901__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06461_ _06460_/Q _06482_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12519__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08200_ _08208_/CLK line[90] VGND VGND VPWR VPWR _08200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05412_ _05424_/CLK line[81] VGND VGND VPWR VPWR _05413_/A sky130_fd_sc_hd__dfxtp_1
X_09180_ _09200_/CLK line[26] VGND VGND VPWR VPWR _09180_/Q sky130_fd_sc_hd__dfxtp_1
X_06392_ _06408_/CLK line[17] VGND VGND VPWR VPWR _06393_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08582__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12816__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08131_ _08131_/A _08162_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05343_ _05342_/Q _05362_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09828__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[2\].TOBUF OVHB\[4\].VALID\[2\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_135_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08062_ _08070_/CLK line[27] VGND VGND VPWR VPWR _08063_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05274_ _05278_/CLK line[18] VGND VGND VPWR VPWR _05275_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07013_ _07012_/Q _07042_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[5\].TOBUF OVHB\[29\].VALID\[5\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06252__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08964_ _08963_/Q _08967_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09563__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07915_ _07915_/CLK _07916_/X VGND VGND VPWR VPWR _07905_/CLK sky130_fd_sc_hd__dlclkp_1
X_08895_ _08895_/CLK _08896_/X VGND VGND VPWR VPWR _08869_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13085__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07846_ _13920_/X wr VGND VGND VPWR VPWR _07846_/X sky130_fd_sc_hd__and2_1
XANTENNA__08179__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08757__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07777_ _13920_/X VGND VGND VPWR VPWR _07777_/Y sky130_fd_sc_hd__inv_2
X_04989_ _04988_/Q _05012_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08476__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06728_ _06740_/CLK line[48] VGND VGND VPWR VPWR _06728_/Q sky130_fd_sc_hd__dfxtp_1
X_09516_ _09515_/Q _09527_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _09427_/CLK line[6] VGND VGND VPWR VPWR _09447_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06659_ _06659_/A _06692_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11333__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06427__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09378_ _09377_/Q _09387_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[5\].VALID\[4\].FF OVHB\[5\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[5\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XMUX.MUX\[14\] _11394_/Z _05584_/Z _13494_/Z _05164_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[14] sky130_fd_sc_hd__mux4_1
X_08329_ _08329_/CLK line[7] VGND VGND VPWR VPWR _08329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09738__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11340_ _11339_/Q _11347_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08642__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11271_ _11251_/CLK line[72] VGND VGND VPWR VPWR _11271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13010_ _13009_/Q _13027_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
X_10222_ _10222_/A _10227_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10153_ _10145_/CLK line[73] VGND VGND VPWR VPWR _10154_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10262__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04939__B2 _04939_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10084_ _10084_/A _10087_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11508__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13912_ _13909_/C _13909_/B _13905_/X _13909_/D VGND VGND VPWR VPWR _06551_/A sky130_fd_sc_hd__and4b_4
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13843_ _13845_/CLK line[110] VGND VGND VPWR VPWR _13843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13723__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[18\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08817__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13774_ _13773_/Q _13797_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_10986_ _10986_/A _10997_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12725_ _12741_/CLK line[111] VGND VGND VPWR VPWR _12725_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11243__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05241__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _12655_/Q _12677_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _11605_/CLK line[97] VGND VGND VPWR VPWR _11608_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _12601_/CLK line[33] VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10437__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08552__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11538_ _11538_/A _11557_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10156__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12074__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11469_ _11479_/CLK line[34] VGND VGND VPWR VPWR _11469_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].V OVHB\[28\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[28\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07168__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13208_ _13207_/Q _13237_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[6\].FF OVHB\[3\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[3\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13139_ _13163_/CLK line[44] VGND VGND VPWR VPWR _13139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09383__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06800__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05961_ _05960_/Q _05992_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11418__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07700_ _07700_/A _07707_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10322__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08680_ _08680_/A _08687_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_05892_ _05902_/CLK line[59] VGND VGND VPWR VPWR _05893_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05416__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07631_ _07633_/CLK line[72] VGND VGND VPWR VPWR _07631_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[7\].TOBUF OVHB\[2\].VALID\[7\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13633__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07562_ _07562_/A _07567_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08727__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06097__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07631__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09301_ _09307_/CLK line[67] VGND VGND VPWR VPWR _09301_/Q sky130_fd_sc_hd__dfxtp_1
X_06513_ _06489_/CLK line[73] VGND VGND VPWR VPWR _06513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12249__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07493_ _07467_/CLK line[9] VGND VGND VPWR VPWR _07493_/Q sky130_fd_sc_hd__dfxtp_1
X_09232_ _09231_/Q _09247_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11731__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06444_ _06443_/Q _06447_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_09163_ _09147_/CLK line[4] VGND VGND VPWR VPWR _09163_/Q sky130_fd_sc_hd__dfxtp_1
X_06375_ _06375_/CLK _06376_/X VGND VGND VPWR VPWR _06353_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09558__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08114_ _08114_/A _08127_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05326_ _13908_/X wr VGND VGND VPWR VPWR _05326_/X sky130_fd_sc_hd__and2_1
XANTENNA__04990__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09094_ _09094_/A _09107_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].CGAND _06551_/A wr VGND VGND VPWR VPWR OVHB\[14\].CGAND/X sky130_fd_sc_hd__and2_4
X_08045_ _08033_/CLK line[5] VGND VGND VPWR VPWR _08045_/Q sky130_fd_sc_hd__dfxtp_1
X_05257_ _13908_/X VGND VGND VPWR VPWR _05257_/Y sky130_fd_sc_hd__inv_2
XOVHB\[31\].VALID\[0\].FF OVHB\[31\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[31\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07078__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].V OVHB\[19\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[19\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05188_ _05214_/CLK line[112] VGND VGND VPWR VPWR _05188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13808__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09996_ _09995_/Q _10017_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09293__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07806__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08947_ _08947_/CLK line[33] VGND VGND VPWR VPWR _08947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10232__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11906__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08878_ _08877_/Q _08897_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07391__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[8\].FF OVHB\[1\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[1\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07829_ _07837_/CLK line[34] VGND VGND VPWR VPWR _07829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10840_ _10840_/A _10857_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07541__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10771_ _10783_/CLK line[99] VGND VGND VPWR VPWR _10771_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12159__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11063__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06157__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _12509_/Q _12537_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_13490_ _13489_/Q _13517_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11998__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12441_ _12449_/CLK line[109] VGND VGND VPWR VPWR _12441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09468__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _12371_/Q _12397_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11323_ _11343_/CLK line[110] VGND VGND VPWR VPWR _11323_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10407__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07566__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11254_ _11253_/Q _11277_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_10205_ _10217_/CLK line[111] VGND VGND VPWR VPWR _10205_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12622__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[11\].FF OVHB\[8\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[8\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11185_ _11191_/CLK line[47] VGND VGND VPWR VPWR _11185_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07716__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10136_ _10136_/A _10157_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11238__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10067_ _10073_/CLK line[33] VGND VGND VPWR VPWR _10068_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09931__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ _13822_/CLK line[88] VGND VGND VPWR VPWR _13827_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[2\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _11345_/CLK sky130_fd_sc_hd__clkbuf_4
X_13757_ _13756_/Q _13762_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10969_ _10977_/CLK line[76] VGND VGND VPWR VPWR _10970_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06067__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ _12708_/CLK line[89] VGND VGND VPWR VPWR _12708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13688_ _13682_/CLK line[25] VGND VGND VPWR VPWR _13688_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12639_ _12638_/Q _12642_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[16\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06160_ _06159_/Q _06167_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08282__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05111_ _05093_/CLK line[72] VGND VGND VPWR VPWR _05112_/A sky130_fd_sc_hd__dfxtp_1
X_06091_ _06077_/CLK line[8] VGND VGND VPWR VPWR _06091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05042_ _05042_/A _05047_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[17\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09850_ _09849_/Q _09877_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06530__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08801_ _08823_/CLK line[109] VGND VGND VPWR VPWR _08801_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[3\].FF OVHB\[28\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[28\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09781_ _09793_/CLK line[45] VGND VGND VPWR VPWR _09782_/A sky130_fd_sc_hd__dfxtp_1
X_06993_ _07001_/CLK line[36] VGND VGND VPWR VPWR _06994_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11148__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05944_ _05943_/Q _05957_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_08732_ _08731_/Q _08757_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05146__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08663_ _08663_/CLK line[46] VGND VGND VPWR VPWR _08664_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10987__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05875_ _05871_/CLK line[37] VGND VGND VPWR VPWR _05875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13363__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07614_ _07613_/Q _07637_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08457__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[10\].VALID\[0\].FF OVHB\[10\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[10\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08594_ _08594_/A _08617_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _07539_/CLK line[47] VGND VGND VPWR VPWR _07545_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[26\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07476_ _07475_/Q _07497_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VOBUF OVHB\[8\].V/Q OVHB\[8\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_06427_ _06421_/CLK line[33] VGND VGND VPWR VPWR _06428_/A sky130_fd_sc_hd__dfxtp_1
X_09215_ _09241_/CLK line[42] VGND VGND VPWR VPWR _09215_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[1\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _08160_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11611__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09146_ _09145_/Q _09177_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06705__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06358_ _06357_/Q _06377_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05309_ _05299_/CLK line[34] VGND VGND VPWR VPWR _05309_/Q sky130_fd_sc_hd__dfxtp_1
X_09077_ _09085_/CLK line[107] VGND VGND VPWR VPWR _09077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06289_ _06285_/CLK line[98] VGND VGND VPWR VPWR _06290_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12292__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08028_ _08027_/Q _08057_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08920__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13538__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09979_ _09978_/Q _09982_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[15\].VALID\[14\].TOBUF OVHB\[15\].VALID\[14\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_12990_ _12990_/CLK _12991_/X VGND VGND VPWR VPWR _12962_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05056__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09106__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10897__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[31\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _11730_/CLK sky130_fd_sc_hd__clkbuf_4
X_11941_ _11872_/A wr VGND VGND VPWR VPWR _11941_/X sky130_fd_sc_hd__and2_1
XANTENNA__13273__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11872_ _11872_/A VGND VGND VPWR VPWR _11872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07271__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[21\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _08860_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[26\].VALID\[5\].FF OVHB\[26\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[26\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13611_ _13610_/Q _13622_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_10823_ _10843_/CLK line[0] VGND VGND VPWR VPWR _10824_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[7\].TOBUF OVHB\[9\].VALID\[7\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12467__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13542_ _13528_/CLK line[86] VGND VGND VPWR VPWR _13542_/Q sky130_fd_sc_hd__dfxtp_1
X_10754_ _10753_/Q _10787_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12186__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13473_ _13472_/Q _13482_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_10685_ _10707_/CLK line[74] VGND VGND VPWR VPWR _10685_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09198__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12424_ _12414_/CLK line[87] VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10137__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ _12355_/A _12362_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[0\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _04975_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08830__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11306_ _11302_/CLK line[88] VGND VGND VPWR VPWR _11306_/Q sky130_fd_sc_hd__dfxtp_1
X_12286_ _12268_/CLK line[24] VGND VGND VPWR VPWR _12287_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13448__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[13\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11237_ _11236_/Q _11242_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12352__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07446__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11168_ _11148_/CLK line[25] VGND VGND VPWR VPWR _11168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10119_ _10118_/Q _10122_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11099_ _11099_/A _11102_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09661__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[25\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13761__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10600__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05660_ _05659_/Q _05677_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_13809_ _13808_/Q _13832_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_05591_ _05575_/CLK line[35] VGND VGND VPWR VPWR _05591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07330_ _07330_/A _07357_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07261_ _07267_/CLK line[45] VGND VGND VPWR VPWR _07261_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[20\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _08475_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__12527__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09000_ _09000_/CLK _09001_/X VGND VGND VPWR VPWR _08972_/CLK sky130_fd_sc_hd__dlclkp_1
X_06212_ _06211_/Q _06237_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[7\].FF OVHB\[24\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[24\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07192_ _07191_/Q _07217_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
X_06143_ _06147_/CLK line[46] VGND VGND VPWR VPWR _06143_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[2\].TOBUF OVHB\[16\].VALID\[2\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_133_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09836__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06074_ _06073_/Q _06097_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[14\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05025_ _05041_/CLK line[47] VGND VGND VPWR VPWR _05025_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12262__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09902_ _09908_/CLK line[86] VGND VGND VPWR VPWR _09902_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13936__A A[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06260__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09833_ _09832_/Q _09842_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09764_ _09760_/CLK line[23] VGND VGND VPWR VPWR _09764_/Q sky130_fd_sc_hd__dfxtp_1
X_06976_ _06975_/Q _07007_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09571__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08715_ _08714_/Q _08722_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_05927_ _05929_/CLK line[75] VGND VGND VPWR VPWR _05927_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13093__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09695_ _09695_/A _09702_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08187__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10510__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05858_ _05857_/Q _05887_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_08646_ _08646_/CLK line[24] VGND VGND VPWR VPWR _08646_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08582_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_05789_ _05799_/CLK line[12] VGND VGND VPWR VPWR _05789_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[7\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _07518_/CLK line[25] VGND VGND VPWR VPWR _07529_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12437__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07459_ _07459_/A _07462_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11341__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09596__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06435__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10470_ _10470_/CLK _10471_/X VGND VGND VPWR VPWR _10466_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09129_ _09128_/Q _09142_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09746__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12140_ _12130_/CLK line[85] VGND VGND VPWR VPWR _12140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13268__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12070_/Q _12082_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[9\].FF OVHB\[22\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[22\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11022_ _11002_/CLK line[86] VGND VGND VPWR VPWR _11023_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06170__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[14\].FF OVHB\[30\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[30\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12900__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[22\].VALID\[1\].TOBUF OVHB\[22\].VALID\[1\].FF/Q OVHB\[22\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].INV _13957_/X VGND VGND VPWR VPWR OVHB\[15\].INV/Y sky130_fd_sc_hd__inv_2
X_12973_ _12972_/Q _12992_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11516__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08097__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11924_ _11934_/CLK line[114] VGND VGND VPWR VPWR _11924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11855_ _11854_/Q _11872_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
X_10806_ _10804_/CLK line[115] VGND VGND VPWR VPWR _10807_/A sky130_fd_sc_hd__dfxtp_1
X_11786_ _11776_/CLK line[51] VGND VGND VPWR VPWR _11786_/Q sky130_fd_sc_hd__dfxtp_1
X_13525_ _13524_/Q _13552_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_10737_ _10736_/Q _10752_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11251__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06345__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13456_ _13468_/CLK line[61] VGND VGND VPWR VPWR _13456_/Q sky130_fd_sc_hd__dfxtp_1
X_10668_ _10656_/CLK line[52] VGND VGND VPWR VPWR _10668_/Q sky130_fd_sc_hd__dfxtp_1
X_12407_ _12406_/Q _12432_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
X_10599_ _10599_/A _10612_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_13387_ _13386_/Q _13412_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08560__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12338_ _12352_/CLK line[62] VGND VGND VPWR VPWR _12339_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13178__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12269_ _12268_/Q _12292_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07176__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11276__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06830_ _06830_/CLK _06831_/X VGND VGND VPWR VPWR _06802_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06761_ _06832_/A wr VGND VGND VPWR VPWR _06761_/X sky130_fd_sc_hd__and2_1
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11426__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08500_ _08480_/CLK line[85] VGND VGND VPWR VPWR _08500_/Q sky130_fd_sc_hd__dfxtp_1
X_05712_ _13909_/X VGND VGND VPWR VPWR _05712_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06692_ _06832_/A VGND VGND VPWR VPWR _06692_/Y sky130_fd_sc_hd__inv_2
X_09480_ _09482_/CLK line[21] VGND VGND VPWR VPWR _09480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05424__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[7\].TOBUF OVHB\[14\].VALID\[7\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08431_ _08431_/A _08442_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_05643_ _05671_/CLK line[64] VGND VGND VPWR VPWR _05643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13641__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08362_ _08358_/CLK line[22] VGND VGND VPWR VPWR _08362_/Q sky130_fd_sc_hd__dfxtp_1
X_05574_ _05573_/Q _05607_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08735__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07313_ _07312_/Q _07322_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
X_08293_ _08292_/Q _08302_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_07244_ _07232_/CLK line[23] VGND VGND VPWR VPWR _07244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07175_ _07174_/Q _07182_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06126_ _06108_/CLK line[24] VGND VGND VPWR VPWR _06126_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[11\].TOBUF OVHB\[9\].VALID\[11\].FF/Q OVHB\[9\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06057_ _06057_/A _06062_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07086__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05008_ _05000_/CLK line[25] VGND VGND VPWR VPWR _05008_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13816__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09816_ _09834_/CLK line[61] VGND VGND VPWR VPWR _09817_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09747_ _09747_/A _09772_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06959_ _06958_/Q _06972_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10240__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09678_ _09694_/CLK line[126] VGND VGND VPWR VPWR _09678_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05334__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08629_ _08628_/Q _08652_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11636_/CLK line[127] VGND VGND VPWR VPWR _11641_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12167__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[2\].VALID\[10\].TOBUF OVHB\[2\].VALID\[10\].FF/Q OVHB\[2\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _11570_/Q _11592_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13308_/CLK line[122] VGND VGND VPWR VPWR _13310_/Q sky130_fd_sc_hd__dfxtp_1
X_10522_ _10520_/CLK line[113] VGND VGND VPWR VPWR _10522_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[6\].TOBUF OVHB\[20\].VALID\[6\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
X_10453_ _10453_/A _10472_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_13241_ _13240_/Q _13272_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09476__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13172_ _13194_/CLK line[59] VGND VGND VPWR VPWR _13172_/Q sky130_fd_sc_hd__dfxtp_1
X_10384_ _10384_/CLK line[50] VGND VGND VPWR VPWR _10384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10415__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12123_ _12123_/A _12152_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05509__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12054_ _12072_/CLK line[60] VGND VGND VPWR VPWR _12054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11005_ _11004_/Q _11032_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12630__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07724__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[13\].CG clk OVHB\[13\].CG/GATE VGND VGND VPWR VPWR OVHB\[13\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_12956_ _12992_/A wr VGND VGND VPWR VPWR _12956_/X sky130_fd_sc_hd__and2_1
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ _11872_/A VGND VGND VPWR VPWR _11907_/Y sky130_fd_sc_hd__inv_2
X_12887_ _12992_/A VGND VGND VPWR VPWR _12887_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11838_ _11846_/CLK line[80] VGND VGND VPWR VPWR _11839_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11769_ _11769_/A _11802_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06075__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13508_ _13507_/Q _13517_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
X_05290_ _05290_/CLK _05291_/X VGND VGND VPWR VPWR _05278_/CLK sky130_fd_sc_hd__dlclkp_1
X_13439_ _13439_/CLK line[39] VGND VGND VPWR VPWR _13439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12805__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08290__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08980_ _08972_/CLK line[63] VGND VGND VPWR VPWR _08980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07931_ _07930_/Q _07952_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12540__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07862_ _07854_/CLK line[49] VGND VGND VPWR VPWR _07863_/A sky130_fd_sc_hd__dfxtp_1
X_09601_ _09600_/Q _09632_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_06813_ _06812_/Q _06832_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07793_ _07792_/Q _07812_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11156__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09532_ _09554_/CLK line[59] VGND VGND VPWR VPWR _09532_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[26\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06744_ _06740_/CLK line[50] VGND VGND VPWR VPWR _06744_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[1\].TOBUF OVHB\[29\].VALID\[1\].FF/Q OVHB\[29\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[18\]_A3 _13605_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09463_ _09462_/Q _09492_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_06675_ _06674_/Q _06692_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13371__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08414_ _08410_/CLK line[60] VGND VGND VPWR VPWR _08414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05626_ _05632_/CLK line[51] VGND VGND VPWR VPWR _05626_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08465__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09394_ _09414_/CLK line[124] VGND VGND VPWR VPWR _09394_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08345_ _08344_/Q _08372_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_05557_ _05556_/Q _05572_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08276_ _08282_/CLK line[125] VGND VGND VPWR VPWR _08276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05488_ _05476_/CLK line[116] VGND VGND VPWR VPWR _05488_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12715__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07227_ _07227_/A _07252_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[12\].TOBUF OVHB\[25\].VALID\[12\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06713__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07158_ _07170_/CLK line[126] VGND VGND VPWR VPWR _07158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06109_ _06108_/Q _06132_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07089_ _07088_/Q _07112_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13546__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12810_ _12810_/A _12817_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_13790_ _13789_/Q _13797_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05064__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05642__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12741_ _12741_/CLK line[104] VGND VGND VPWR VPWR _12741_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].CG clk OVHB\[8\].CGAND/X VGND VGND VPWR VPWR OVHB\[8\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13281__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05999__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05361__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08375__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12672_/A _12677_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[0\]_A1 _10894_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11605_/CLK line[105] VGND VGND VPWR VPWR _11623_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _11553_/Q _11557_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _10505_/CLK _10506_/X VGND VGND VPWR VPWR _10473_/CLK sky130_fd_sc_hd__dlclkp_1
X_11485_ _11485_/CLK _11486_/X VGND VGND VPWR VPWR _11479_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_100_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06623__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13224_ _13223_/Q _13237_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_10436_ _13931_/X wr VGND VGND VPWR VPWR _10436_/X sky130_fd_sc_hd__and2_1
XFILLER_128_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10145__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13155_ _13163_/CLK line[37] VGND VGND VPWR VPWR _13155_/Q sky130_fd_sc_hd__dfxtp_1
X_10367_ _13931_/X VGND VGND VPWR VPWR _10367_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05239__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05817__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12106_ _12105_/Q _12117_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_13086_ _13086_/A _13097_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_10298_ _10314_/CLK line[16] VGND VGND VPWR VPWR _10298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13456__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12037_ _12019_/CLK line[38] VGND VGND VPWR VPWR _12037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05536__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07454__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13988_ _13990_/B _13990_/A _13982_/X _13990_/D VGND VGND VPWR VPWR _13988_/X sky130_fd_sc_hd__and4b_4
XFILLER_46_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12939_ _12937_/CLK line[66] VGND VGND VPWR VPWR _12939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11704__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06460_ _06464_/CLK line[63] VGND VGND VPWR VPWR _06460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05702__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05411_ _05410_/Q _05432_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
X_06391_ _06391_/A _06412_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08130_ _08134_/CLK line[58] VGND VGND VPWR VPWR _08131_/A sky130_fd_sc_hd__dfxtp_1
X_05342_ _05332_/CLK line[49] VGND VGND VPWR VPWR _05342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04934__A2_N _04934_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08061_ _08060_/Q _08092_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_05273_ _05272_/Q _05292_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[3\].TOBUF OVHB\[2\].VALID\[3\].FF/Q OVHB\[2\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_105_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07012_ _07030_/CLK line[59] VGND VGND VPWR VPWR _07012_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07629__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[6\].TOBUF OVHB\[27\].VALID\[6\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__10055__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08963_ _08947_/CLK line[41] VGND VGND VPWR VPWR _08963_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12270__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07914_ _07913_/Q _07917_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04988__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08894_ _08894_/A _08897_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07364__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07845_ _07845_/CLK _07846_/X VGND VGND VPWR VPWR _07837_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_57_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[10\].CGAND _13908_/X wr VGND VGND VPWR VPWR OVHB\[10\].CGAND/X sky130_fd_sc_hd__and2_4
X_07776_ _13920_/X wr VGND VGND VPWR VPWR _07776_/X sky130_fd_sc_hd__and2_1
X_04988_ _05000_/CLK line[30] VGND VGND VPWR VPWR _04988_/Q sky130_fd_sc_hd__dfxtp_1
X_09515_ _09507_/CLK line[37] VGND VGND VPWR VPWR _09515_/Q sky130_fd_sc_hd__dfxtp_1
X_06727_ _06832_/A VGND VGND VPWR VPWR _06727_/Y sky130_fd_sc_hd__inv_2
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09446_ _09445_/Q _09457_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06658_ _06682_/CLK line[16] VGND VGND VPWR VPWR _06659_/A sky130_fd_sc_hd__dfxtp_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05612__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[31\]_A0 _10871_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05609_ _05608_/Q _05642_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_09377_ _09365_/CLK line[102] VGND VGND VPWR VPWR _09377_/Q sky130_fd_sc_hd__dfxtp_1
X_06589_ _06588_/Q _06622_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08328_ _08327_/Q _08337_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12445__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08259_ _08257_/CLK line[103] VGND VGND VPWR VPWR _08259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07539__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06443__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11270_ _11269_/Q _11277_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[8\].VALID\[9\].FF OVHB\[8\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[8\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10221_ _10217_/CLK line[104] VGND VGND VPWR VPWR _10222_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09754__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10152_ _10151_/Q _10157_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_10083_ _10073_/CLK line[41] VGND VGND VPWR VPWR _10084_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ _13909_/B _13909_/C _13905_/X _13909_/D VGND VGND VPWR VPWR _06272_/A sky130_fd_sc_hd__and4b_4
X_13842_ _13842_/A _13867_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13773_ _13763_/CLK line[78] VGND VGND VPWR VPWR _13773_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[24\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10985_ _10977_/CLK line[69] VGND VGND VPWR VPWR _10986_/A sky130_fd_sc_hd__dfxtp_1
X_12724_ _12723_/Q _12747_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06618__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12655_ _12667_/CLK line[79] VGND VGND VPWR VPWR _12655_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _11606_/A _11627_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[8\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[12\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12586_ _12585_/Q _12607_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _11535_/CLK line[65] VGND VGND VPWR VPWR _11538_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06353__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11468_ _11467_/Q _11487_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_13207_ _13213_/CLK line[75] VGND VGND VPWR VPWR _13207_/Q sky130_fd_sc_hd__dfxtp_1
X_10419_ _10405_/CLK line[66] VGND VGND VPWR VPWR _10419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[24\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11399_ _11395_/CLK line[2] VGND VGND VPWR VPWR _11400_/A sky130_fd_sc_hd__dfxtp_1
X_13138_ _13138_/A _13167_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13186__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13069_ _13075_/CLK line[12] VGND VGND VPWR VPWR _13069_/Q sky130_fd_sc_hd__dfxtp_1
X_05960_ _05984_/CLK line[90] VGND VGND VPWR VPWR _05960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05891_ _05891_/A _05922_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07630_ _07629_/Q _07637_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[8\].TOBUF OVHB\[0\].VALID\[8\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07561_ _07539_/CLK line[40] VGND VGND VPWR VPWR _07562_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11434__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ _09299_/Q _09317_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_06512_ _06512_/A _06517_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06528__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07492_ _07491_/Q _07497_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09231_ _09241_/CLK line[35] VGND VGND VPWR VPWR _09231_/Q sky130_fd_sc_hd__dfxtp_1
X_06443_ _06421_/CLK line[41] VGND VGND VPWR VPWR _06443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11731__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08743__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06374_ _06373_/Q _06377_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_09162_ _09161_/Q _09177_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_08113_ _08113_/CLK line[36] VGND VGND VPWR VPWR _08114_/A sky130_fd_sc_hd__dfxtp_1
X_05325_ _05325_/CLK _05326_/X VGND VGND VPWR VPWR _05299_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09093_ _09085_/CLK line[100] VGND VGND VPWR VPWR _09094_/A sky130_fd_sc_hd__dfxtp_1
X_08044_ _08044_/A _08057_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_05256_ _13908_/X wr VGND VGND VPWR VPWR _05256_/X sky130_fd_sc_hd__and2_1
X_05187_ _05152_/A VGND VGND VPWR VPWR _05187_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[17\].VALID\[1\].FF OVHB\[17\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[17\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09995_ _10011_/CLK line[15] VGND VGND VPWR VPWR _09995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11609__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08946_ _08945_/Q _08967_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VOBUF OVHB\[4\].V/Q OVHB\[4\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
XANTENNA__07094__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07672__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11906__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08877_ _08869_/CLK line[1] VGND VGND VPWR VPWR _08877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13824__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07391__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07828_ _07827_/Q _07847_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08918__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07759_ _07773_/CLK line[2] VGND VGND VPWR VPWR _07759_/Q sky130_fd_sc_hd__dfxtp_1
X_10770_ _10770_/A _10787_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05342__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09429_ _09427_/CLK line[12] VGND VGND VPWR VPWR _09429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12440_ _12439_/Q _12467_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08653__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[10\].TOBUF OVHB\[15\].VALID\[10\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12175__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _12387_/CLK line[77] VGND VGND VPWR VPWR _12371_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07269__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07847__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11322_ _11321_/Q _11347_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07566__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11253_ _11251_/CLK line[78] VGND VGND VPWR VPWR _11253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09484__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[3\].TOBUF OVHB\[9\].VALID\[3\].FF/Q OVHB\[9\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XFILLER_122_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10204_ _10203_/Q _10227_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11184_ _11183_/Q _11207_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10423__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10135_ _10145_/CLK line[79] VGND VGND VPWR VPWR _10136_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05517__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10066_ _10065_/Q _10087_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13734__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08828__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[3\].FF OVHB\[15\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[15\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07732__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13825_ _13824_/Q _13832_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13756_ _13746_/CLK line[56] VGND VGND VPWR VPWR _13756_/Q sky130_fd_sc_hd__dfxtp_1
X_10968_ _10967_/Q _10997_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
X_12707_ _12706_/Q _12712_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[12\].FF OVHB\[31\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[31\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13687_ _13686_/Q _13692_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_10899_ _10903_/CLK line[44] VGND VGND VPWR VPWR _10899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09659__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ _12638_/CLK line[57] VGND VGND VPWR VPWR _12638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[22\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12085__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12569_ _12569_/A _12572_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05110_ _05109_/Q _05117_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06083__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06090_ _06090_/A _06097_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05041_ _05041_/CLK line[40] VGND VGND VPWR VPWR _05042_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12813__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07907__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09394__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08800_ _08800_/A _08827_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10333__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09780_ _09780_/A _09807_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06992_ _06992_/A _07007_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__04919__A1_N A_h[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08731_ _08749_/CLK line[77] VGND VGND VPWR VPWR _08731_/Q sky130_fd_sc_hd__dfxtp_1
X_05943_ _05929_/CLK line[68] VGND VGND VPWR VPWR _05943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[14\].FF OVHB\[21\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[21\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08662_ _08661_/Q _08687_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_05874_ _05873_/Q _05887_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07642__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07613_ _07633_/CLK line[78] VGND VGND VPWR VPWR _07613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ _08609_/CLK line[14] VGND VGND VPWR VPWR _08594_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11164__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07544_ _07544_/A _07567_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06258__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09212__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ _07467_/CLK line[15] VGND VGND VPWR VPWR _07475_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09569__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09214_ _09213_/Q _09247_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
X_06426_ _06426_/A _06447_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08473__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[5\].FF OVHB\[13\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[13\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09145_ _09147_/CLK line[10] VGND VGND VPWR VPWR _09145_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10508__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[9\].FF OVHB\[30\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[30\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06357_ _06353_/CLK line[1] VGND VGND VPWR VPWR _06357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05308_ _05308_/A _05327_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_06288_ _06287_/Q _06307_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
X_09076_ _09075_/Q _09107_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12723__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08027_ _08033_/CLK line[11] VGND VGND VPWR VPWR _08027_/Q sky130_fd_sc_hd__dfxtp_1
X_05239_ _05253_/CLK line[2] VGND VGND VPWR VPWR _05239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07817__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05187__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06721__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11339__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10821__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09978_ _09978_/CLK line[121] VGND VGND VPWR VPWR _09978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08929_ _08928_/Q _08932_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11940_ _11940_/CLK _11941_/X VGND VGND VPWR VPWR _11934_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08648__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09106__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11871_ _11872_/A wr VGND VGND VPWR VPWR _11871_/X sky130_fd_sc_hd__and2_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11074__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13610_ _13598_/CLK line[117] VGND VGND VPWR VPWR _13610_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06168__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10822_ _13932_/X VGND VGND VPWR VPWR _10822_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05072__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[8\].TOBUF OVHB\[7\].VALID\[8\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_13541_ _13540_/Q _13552_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_10753_ _10783_/CLK line[96] VGND VGND VPWR VPWR _10753_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DECH.DEC0.AND2_B A_h[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08383__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13472_ _13468_/CLK line[54] VGND VGND VPWR VPWR _13472_/Q sky130_fd_sc_hd__dfxtp_1
X_10684_ _10683_/Q _10717_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12423_ _12422_/Q _12432_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_12354_ _12352_/CLK line[55] VGND VGND VPWR VPWR _12355_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06481__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11305_ _11304_/Q _11312_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_12285_ _12284_/Q _12292_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[7\].FF OVHB\[11\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[11\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06631__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11236_ _11216_/CLK line[56] VGND VGND VPWR VPWR _11236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11249__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10153__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11167_ _11166_/Q _11172_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05247__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10118_ _10100_/CLK line[57] VGND VGND VPWR VPWR _10118_/Q sky130_fd_sc_hd__dfxtp_1
X_11098_ _11090_/CLK line[121] VGND VGND VPWR VPWR _11099_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13464__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08558__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10049_ _10048_/Q _10052_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13761__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05590_ _05589_/Q _05607_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_13808_ _13822_/CLK line[94] VGND VGND VPWR VPWR _13808_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06656__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13739_ _13738_/Q _13762_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11712__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06806__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07260_ _07259_/Q _07287_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_06211_ _06223_/CLK line[77] VGND VGND VPWR VPWR _06211_/Q sky130_fd_sc_hd__dfxtp_1
X_07191_ _07183_/CLK line[13] VGND VGND VPWR VPWR _07191_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10328__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06142_ _06141_/Q _06167_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[19\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _07845_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13639__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[14\].VALID\[3\].TOBUF OVHB\[14\].VALID\[3\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_06073_ _06077_/CLK line[14] VGND VGND VPWR VPWR _06073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05024_ _05023_/Q _05047_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_09901_ _09901_/A _09912_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XDEC.DEC0.AND0 A[7] A[8] VGND VGND VPWR VPWR _13944_/D sky130_fd_sc_hd__nor2_2
XFILLER_99_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10063__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09832_ _09834_/CLK line[54] VGND VGND VPWR VPWR _09832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05157__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10998__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09763_ _09762_/Q _09772_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_06975_ _07001_/CLK line[42] VGND VGND VPWR VPWR _06975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08714_ _08710_/CLK line[55] VGND VGND VPWR VPWR _08714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04996__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05926_ _05925_/Q _05957_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
X_09694_ _09694_/CLK line[119] VGND VGND VPWR VPWR _09695_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07372__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08645_ _08644_/Q _08652_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_05857_ _05871_/CLK line[43] VGND VGND VPWR VPWR _05857_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _08560_/CLK line[120] VGND VGND VPWR VPWR _08577_/A sky130_fd_sc_hd__dfxtp_1
X_05788_ _05788_/A _05817_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[21\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07527_ _07526_/Q _07532_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09299__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09877__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ _07446_/CLK line[121] VGND VGND VPWR VPWR _07459_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05620__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06409_ _06409_/A _06412_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09596__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07389_ _07388_/Q _07392_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[14\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09128_ _09116_/CLK line[116] VGND VGND VPWR VPWR _09128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12453__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09059_ _09058_/Q _09072_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07547__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12070_ _12072_/CLK line[53] VGND VGND VPWR VPWR _12070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11021_ _11020_/Q _11032_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09762__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08021__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10701__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12972_ _12962_/CLK line[81] VGND VGND VPWR VPWR _12972_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[2\].TOBUF OVHB\[20\].VALID\[2\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_100_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11923_ _11923_/A _11942_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11382__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11854_ _11846_/CLK line[82] VGND VGND VPWR VPWR _11854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10805_ _10804_/Q _10822_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04920__B1 A_h[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12628__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11785_ _11785_/A _11802_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_13524_ _13528_/CLK line[92] VGND VGND VPWR VPWR _13524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10736_ _10728_/CLK line[83] VGND VGND VPWR VPWR _10736_/Q sky130_fd_sc_hd__dfxtp_1
X_13455_ _13454_/Q _13482_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10667_ _10667_/A _10682_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09937__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12406_ _12414_/CLK line[93] VGND VGND VPWR VPWR _12406_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13386_ _13394_/CLK line[29] VGND VGND VPWR VPWR _13386_/Q sky130_fd_sc_hd__dfxtp_1
X_10598_ _10594_/CLK line[20] VGND VGND VPWR VPWR _10599_/A sky130_fd_sc_hd__dfxtp_1
X_12337_ _12336_/Q _12362_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12363__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06361__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12268_ _12268_/CLK line[30] VGND VGND VPWR VPWR _12268_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[0\].FF OVHB\[4\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[4\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[25\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11219_ _11218_/Q _11242_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[15\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11557__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12199_ _12199_/A _12222_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09672__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11276__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13194__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06760_ _06760_/CLK _06761_/X VGND VGND VPWR VPWR _06740_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08288__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05711_ _13909_/X wr VGND VGND VPWR VPWR _05711_/X sky130_fd_sc_hd__and2_1
X_06691_ _06832_/A wr VGND VGND VPWR VPWR _06691_/X sky130_fd_sc_hd__and2_1
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08430_ _08410_/CLK line[53] VGND VGND VPWR VPWR _08431_/A sky130_fd_sc_hd__dfxtp_1
X_05642_ _13909_/X VGND VGND VPWR VPWR _05642_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[8\].TOBUF OVHB\[12\].VALID\[8\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07920__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08361_ _08361_/A _08372_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12538__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05573_ _05575_/CLK line[32] VGND VGND VPWR VPWR _05573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11442__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07312_ _07292_/CLK line[54] VGND VGND VPWR VPWR _07312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06536__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08292_ _08282_/CLK line[118] VGND VGND VPWR VPWR _08292_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[12\].TOBUF OVHB\[5\].VALID\[12\].FF/Q OVHB\[5\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_20_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[8\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07243_ _07242_/Q _07252_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09847__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08751__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07174_ _07170_/CLK line[119] VGND VGND VPWR VPWR _07174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13369__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13947__A A_h[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06125_ _06125_/A _06132_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12851__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06056_ _06050_/CLK line[120] VGND VGND VPWR VPWR _06057_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05007_ _05006_/Q _05012_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09815_ _09814_/Q _09842_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11617__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08198__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09746_ _09760_/CLK line[29] VGND VGND VPWR VPWR _09747_/A sky130_fd_sc_hd__dfxtp_1
X_06958_ _06960_/CLK line[20] VGND VGND VPWR VPWR _06958_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[2\].FF OVHB\[2\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[2\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05909_ _05909_/A _05922_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_09677_ _09677_/A _09702_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_06889_ _06888_/Q _06902_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08646_/CLK line[30] VGND VGND VPWR VPWR _08628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08926__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08559_/A _08582_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11352__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _11588_/CLK line[95] VGND VGND VPWR VPWR _11570_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05350__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10521_ _10521_/A _10542_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08661__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13240_ _13254_/CLK line[90] VGND VGND VPWR VPWR _13240_/Q sky130_fd_sc_hd__dfxtp_1
X_10452_ _10466_/CLK line[81] VGND VGND VPWR VPWR _10453_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13279__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12183__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13171_ _13170_/Q _13202_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_10383_ _10382_/Q _10402_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07277__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[16\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12122_ _12130_/CLK line[91] VGND VGND VPWR VPWR _12123_/A sky130_fd_sc_hd__dfxtp_1
X_12053_ _12052_/Q _12082_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11004_ _11002_/CLK line[92] VGND VGND VPWR VPWR _11004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11527__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10431__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08686__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05525__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12955_ _12955_/CLK _12956_/X VGND VGND VPWR VPWR _12937_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13742__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11906_ _11872_/A wr VGND VGND VPWR VPWR _11906_/X sky130_fd_sc_hd__and2_1
XANTENNA__08836__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12886_ _12992_/A wr VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__and2_1
XANTENNA__12358__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11837_ _11872_/A VGND VGND VPWR VPWR _11837_/Y sky130_fd_sc_hd__inv_2
XMUX.MUX\[1\] _04958_/Z _13428_/Z _13498_/Z _13568_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[1] sky130_fd_sc_hd__mux4_1
XFILLER_53_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11768_ _11776_/CLK line[48] VGND VGND VPWR VPWR _11769_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05260__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[4\].FF OVHB\[0\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[0\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _13497_/CLK line[70] VGND VGND VPWR VPWR _13507_/Q sky130_fd_sc_hd__dfxtp_1
X_10719_ _10718_/Q _10752_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_11699_ _11698_/Q _11732_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
X_13438_ _13437_/Q _13447_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[14\].TOBUF OVHB\[28\].VALID\[14\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__12093__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10606__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13369_ _13347_/CLK line[7] VGND VGND VPWR VPWR _13370_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07187__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06091__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[26\].VALID\[14\].FF OVHB\[26\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[26\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07930_ _07946_/CLK line[95] VGND VGND VPWR VPWR _07930_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10191__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07861_ _07860_/Q _07882_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
X_09600_ _09626_/CLK line[90] VGND VGND VPWR VPWR _09600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10341__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06812_ _06802_/CLK line[81] VGND VGND VPWR VPWR _06812_/Q sky130_fd_sc_hd__dfxtp_1
X_07792_ _07788_/CLK line[17] VGND VGND VPWR VPWR _07792_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05435__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09531_ _09530_/Q _09562_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_06743_ _06742_/Q _06762_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[26\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[13\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09462_ _09482_/CLK line[27] VGND VGND VPWR VPWR _09462_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[2\].TOBUF OVHB\[27\].VALID\[2\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06674_ _06682_/CLK line[18] VGND VGND VPWR VPWR _06674_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07650__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08413_ _08412_/Q _08442_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05625_ _05624_/Q _05642_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12268__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09393_ _09392_/Q _09422_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[13\].TOBUF OVHB\[21\].VALID\[13\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ _08358_/CLK line[28] VGND VGND VPWR VPWR _08344_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06266__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05556_ _05568_/CLK line[19] VGND VGND VPWR VPWR _05556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08275_ _08274_/Q _08302_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10366__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05487_ _05487_/A _05502_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09577__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07226_ _07232_/CLK line[29] VGND VGND VPWR VPWR _07227_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].INV _13956_/X VGND VGND VPWR VPWR OVHB\[14\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_4_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10516__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07157_ _07156_/Q _07182_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[6\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06108_ _06108_/CLK line[30] VGND VGND VPWR VPWR _06108_/Q sky130_fd_sc_hd__dfxtp_1
X_07088_ _07098_/CLK line[94] VGND VGND VPWR VPWR _07088_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].INV _13977_/X VGND VGND VPWR VPWR OVHB\[29\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__12731__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06039_ _06038_/Q _06062_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07825__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09729_ _09721_/CLK line[7] VGND VGND VPWR VPWR _09730_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12740_ _12739_/Q _12747_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12667_/CLK line[72] VGND VGND VPWR VPWR _12672_/A sky130_fd_sc_hd__dfxtp_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11082__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06176__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11621_/Q _11627_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[0\]_A2 _05084_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[19\].VALID\[8\].TOBUF OVHB\[19\].VALID\[8\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12906__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _11535_/CLK line[73] VGND VGND VPWR VPWR _11553_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08391__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10504_ _10504_/A _10507_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11484_ _11483_/Q _11487_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13223_ _13213_/CLK line[68] VGND VGND VPWR VPWR _13223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13587__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10435_ _10435_/CLK _10436_/X VGND VGND VPWR VPWR _10405_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[23\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13154_ _13153_/Q _13167_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10366_ _13931_/X wr VGND VGND VPWR VPWR _10366_/X sky130_fd_sc_hd__and2_1
XDATA\[9\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _13760_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12105_ _12109_/CLK line[69] VGND VGND VPWR VPWR _12105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13085_ _13075_/CLK line[5] VGND VGND VPWR VPWR _13086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10297_ _13931_/X VGND VGND VPWR VPWR _10297_/Y sky130_fd_sc_hd__inv_2
X_12036_ _12035_/Q _12047_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11257__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09950__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ _13990_/A _13990_/B _13982_/X _13990_/D VGND VGND VPWR VPWR _13987_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__13472__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08566__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12938_ _12937_/Q _12957_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12869_ _12881_/CLK line[34] VGND VGND VPWR VPWR _12869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[23\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05410_ _05424_/CLK line[95] VGND VGND VPWR VPWR _05410_/Q sky130_fd_sc_hd__dfxtp_1
X_06390_ _06408_/CLK line[31] VGND VGND VPWR VPWR _06391_/A sky130_fd_sc_hd__dfxtp_1
X_05341_ _05341_/A _05362_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11720__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[29\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _11100_/CLK sky130_fd_sc_hd__clkbuf_4
X_08060_ _08070_/CLK line[26] VGND VGND VPWR VPWR _08060_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06814__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05272_ _05278_/CLK line[17] VGND VGND VPWR VPWR _05272_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[1\].FF OVHB\[25\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[25\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07011_ _07010_/Q _07042_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[4\].TOBUF OVHB\[0\].VALID\[4\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[25\].VALID\[7\].TOBUF OVHB\[25\].VALID\[7\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13647__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08962_ _08961_/Q _08967_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07913_ _07905_/CLK line[73] VGND VGND VPWR VPWR _07913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08893_ _08869_/CLK line[9] VGND VGND VPWR VPWR _08894_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[8\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _13375_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10071__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07844_ _07843_/Q _07847_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05165__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07775_ _07775_/CLK _07776_/X VGND VGND VPWR VPWR _07773_/CLK sky130_fd_sc_hd__dlclkp_1
X_04987_ _04987_/A _05012_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13382__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13960__A A_h[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09514_ _09513_/Q _09527_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06726_ _06832_/A wr VGND VGND VPWR VPWR _06726_/X sky130_fd_sc_hd__and2_1
XANTENNA__07380__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09445_ _09427_/CLK line[5] VGND VGND VPWR VPWR _09445_/Q sky130_fd_sc_hd__dfxtp_1
X_06657_ _06832_/A VGND VGND VPWR VPWR _06657_/Y sky130_fd_sc_hd__inv_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05608_ _05632_/CLK line[48] VGND VGND VPWR VPWR _05608_/Q sky130_fd_sc_hd__dfxtp_1
X_09376_ _09375_/Q _09387_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[31\]_A1 _13461_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06588_ _06596_/CLK line[112] VGND VGND VPWR VPWR _06588_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VOBUF OVHB\[0\].V/Q OVHB\[0\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_08327_ _08329_/CLK line[6] VGND VGND VPWR VPWR _08327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[11\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05539_ _05538_/Q _05572_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[12\].FF OVHB\[22\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[22\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11630__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08258_ _08258_/A _08267_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_07209_ _07183_/CLK line[7] VGND VGND VPWR VPWR _07209_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10246__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08189_ _08175_/CLK line[71] VGND VGND VPWR VPWR _08189_/Q sky130_fd_sc_hd__dfxtp_1
X_10220_ _10220_/A _10227_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[28\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _10715_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[4\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13557__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12461__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10151_ _10145_/CLK line[72] VGND VGND VPWR VPWR _10151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[3\].FF OVHB\[23\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[23\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07555__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10082_ _10082_/A _10087_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13910_ _13909_/C _13909_/B _13905_/X _13909_/D VGND VGND VPWR VPWR _13910_/X sky130_fd_sc_hd__and4bb_4
XANTENNA_DATA\[4\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13841_ _13845_/CLK line[109] VGND VGND VPWR VPWR _13842_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11805__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[14\].FF OVHB\[12\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[12\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[6\].TOBUF OVHB\[31\].VALID\[6\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13772_ _13771_/Q _13797_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07290__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10984_ _10983_/Q _10997_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05803__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[30\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12723_ _12741_/CLK line[110] VGND VGND VPWR VPWR _12723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _12653_/Q _12677_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11605_/CLK line[111] VGND VGND VPWR VPWR _11606_/A sky130_fd_sc_hd__dfxtp_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12601_/CLK line[47] VGND VGND VPWR VPWR _12585_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.MUX\[8\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ _11535_/Q _11557_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ _11479_/CLK line[33] VGND VGND VPWR VPWR _11467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_MUX.MUX\[16\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13206_ _13205_/Q _13237_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10418_ _10418_/A _10437_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
X_11398_ _11397_/Q _11417_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_13137_ _13163_/CLK line[43] VGND VGND VPWR VPWR _13138_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12371__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10349_ _10341_/CLK line[34] VGND VGND VPWR VPWR _10349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07465__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13068_ _13067_/Q _13097_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[27\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _10330_/CLK sky130_fd_sc_hd__clkbuf_4
X_12019_ _12019_/CLK line[44] VGND VGND VPWR VPWR _12019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05890_ _05902_/CLK line[58] VGND VGND VPWR VPWR _05891_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09680__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _07460_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[5\].FF OVHB\[21\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[21\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07560_ _07559_/Q _07567_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08296__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05713__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06511_ _06489_/CLK line[72] VGND VGND VPWR VPWR _06512_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07491_ _07467_/CLK line[8] VGND VGND VPWR VPWR _07491_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12396__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09230_ _09229_/Q _09247_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_06442_ _06441_/Q _06447_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09161_ _09147_/CLK line[3] VGND VGND VPWR VPWR _09161_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12546__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06373_ _06353_/CLK line[9] VGND VGND VPWR VPWR _06373_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].CG clk OVHB\[26\].CGAND/X VGND VGND VPWR VPWR OVHB\[26\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_08112_ _08112_/A _08127_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06544__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05324_ _05324_/A _05327_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_09092_ _09091_/Q _09107_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[12\].TOBUF OVHB\[18\].VALID\[12\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08043_ _08033_/CLK line[4] VGND VGND VPWR VPWR _08044_/A sky130_fd_sc_hd__dfxtp_1
X_05255_ _05255_/CLK _05256_/X VGND VGND VPWR VPWR _05253_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_31_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09855__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05186_ _05152_/A wr VGND VGND VPWR VPWR _05186_/X sky130_fd_sc_hd__and2_1
XFILLER_115_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _09993_/Q _10017_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08945_ _08947_/CLK line[47] VGND VGND VPWR VPWR _08945_/Q sky130_fd_sc_hd__dfxtp_1
X_08876_ _08875_/Q _08897_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
X_07827_ _07837_/CLK line[33] VGND VGND VPWR VPWR _07827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[29\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06719__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07758_ _07757_/Q _07777_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[11\].TOBUF OVHB\[11\].VALID\[11\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_06709_ _06711_/CLK line[34] VGND VGND VPWR VPWR _06709_/Q sky130_fd_sc_hd__dfxtp_1
X_07689_ _07679_/CLK line[98] VGND VGND VPWR VPWR _07689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[16\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _07075_/CLK sky130_fd_sc_hd__clkbuf_4
X_09428_ _09428_/A _09457_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].CGAND _13272_/A wr VGND VGND VPWR VPWR OVHB\[7\].CGAND/X sky130_fd_sc_hd__and2_4
X_09359_ _09365_/CLK line[108] VGND VGND VPWR VPWR _09360_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11360__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06454__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12370_ _12369_/Q _12397_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11321_ _11343_/CLK line[109] VGND VGND VPWR VPWR _11321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11252_ _11251_/Q _11277_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13287__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10203_ _10217_/CLK line[110] VGND VGND VPWR VPWR _10203_/Q sky130_fd_sc_hd__dfxtp_1
X_11183_ _11191_/CLK line[46] VGND VGND VPWR VPWR _11183_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[4\].TOBUF OVHB\[7\].VALID\[4\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_79_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10134_ _10134_/A _10157_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10065_ _10073_/CLK line[47] VGND VGND VPWR VPWR _10065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__04933__A2_N _04933_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11535__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06629__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13824_ _13822_/CLK line[87] VGND VGND VPWR VPWR _13824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05533__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09005__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13755_ _13754_/Q _13762_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
X_10967_ _10977_/CLK line[75] VGND VGND VPWR VPWR _10967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13750__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[2\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08844__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12706_ _12708_/CLK line[88] VGND VGND VPWR VPWR _12706_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ _10897_/Q _10927_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
X_13686_ _13682_/CLK line[24] VGND VGND VPWR VPWR _13686_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[8\].FF OVHB\[18\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[18\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _12636_/Q _12642_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[15\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _06690_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_129_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12568_ _12560_/CLK line[25] VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11519_ _11518_/Q _11522_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_12499_ _12498_/Q _12502_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05040_ _05039_/Q _05047_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07195__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05708__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06991_ _07001_/CLK line[35] VGND VGND VPWR VPWR _06992_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[31\].VALID\[11\].TOBUF OVHB\[31\].VALID\[11\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[21\]_A0 _10881_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08730_ _08729_/Q _08757_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_05942_ _05941_/Q _05957_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08661_ _08663_/CLK line[45] VGND VGND VPWR VPWR _08661_/Q sky130_fd_sc_hd__dfxtp_1
X_05873_ _05871_/CLK line[36] VGND VGND VPWR VPWR _05873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07612_ _07611_/Q _07637_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08592_ _08591_/Q _08617_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05443__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07543_ _07539_/CLK line[46] VGND VGND VPWR VPWR _07544_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13660__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07474_ _07473_/Q _07497_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09213_ _09241_/CLK line[32] VGND VGND VPWR VPWR _09213_/Q sky130_fd_sc_hd__dfxtp_1
X_06425_ _06421_/CLK line[47] VGND VGND VPWR VPWR _06426_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12276__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09144_ _09143_/Q _09177_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_06356_ _06356_/A _06377_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05307_ _05299_/CLK line[33] VGND VGND VPWR VPWR _05308_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09075_ _09085_/CLK line[106] VGND VGND VPWR VPWR _09075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06287_ _06285_/CLK line[97] VGND VGND VPWR VPWR _06287_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09585__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08026_ _08025_/Q _08057_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_05238_ _05238_/A _05257_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10524__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05169_ _05157_/CLK line[98] VGND VGND VPWR VPWR _05170_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_115_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05618__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09977_ _09977_/A _09982_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13835__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10821__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08928_ _08922_/CLK line[25] VGND VGND VPWR VPWR _08928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07833__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08859_ _08859_/A _08862_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11870_ _11870_/CLK _11871_/X VGND VGND VPWR VPWR _11846_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10821_ _13932_/X wr VGND VGND VPWR VPWR _10821_/X sky130_fd_sc_hd__and2_1
XFILLER_26_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13540_ _13528_/CLK line[85] VGND VGND VPWR VPWR _13540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10752_ _13932_/X VGND VGND VPWR VPWR _10752_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[9\].TOBUF OVHB\[5\].VALID\[9\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[3\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13471_ _13470_/Q _13482_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_10683_ _10707_/CLK line[64] VGND VGND VPWR VPWR _10683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11090__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06184__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12422_ _12414_/CLK line[86] VGND VGND VPWR VPWR _12422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06762__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12353_ _12352_/Q _12362_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12914__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[23\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06481__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09495__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11304_ _11302_/CLK line[87] VGND VGND VPWR VPWR _11304_/Q sky130_fd_sc_hd__dfxtp_1
X_12284_ _12268_/CLK line[23] VGND VGND VPWR VPWR _12284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11235_ _11235_/A _11242_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11166_ _11148_/CLK line[24] VGND VGND VPWR VPWR _11166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10117_ _10116_/Q _10122_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11097_ _11096_/Q _11102_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07743__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[14\].FF OVHB\[3\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[3\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10048_ _10042_/CLK line[25] VGND VGND VPWR VPWR _10048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11265__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06359__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06937__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13807_ _13806_/Q _13832_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06656__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11999_ _11998_/Q _12012_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08574__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13738_ _13746_/CLK line[62] VGND VGND VPWR VPWR _13738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13669_ _13669_/A _13692_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06210_ _06209_/Q _06237_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
X_07190_ _07190_/A _07217_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06141_ _06147_/CLK line[45] VGND VGND VPWR VPWR _06141_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].V OVHB\[4\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[4\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12824__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07918__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06822__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06072_ _06071_/Q _06097_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[4\].TOBUF OVHB\[12\].VALID\[4\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_05023_ _05041_/CLK line[46] VGND VGND VPWR VPWR _05023_/Q sky130_fd_sc_hd__dfxtp_1
X_09900_ _09908_/CLK line[85] VGND VGND VPWR VPWR _09901_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDEC.DEC0.AND1 A[8] A[7] VGND VGND VPWR VPWR _13909_/D sky130_fd_sc_hd__and2b_2
X_09831_ _09830_/Q _09842_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_06974_ _06973_/Q _07007_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08749__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09762_ _09760_/CLK line[22] VGND VGND VPWR VPWR _09762_/Q sky130_fd_sc_hd__dfxtp_1
X_08713_ _08712_/Q _08722_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05925_ _05929_/CLK line[74] VGND VGND VPWR VPWR _05925_/Q sky130_fd_sc_hd__dfxtp_1
X_09693_ _09692_/Q _09702_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11175__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08644_ _08646_/CLK line[23] VGND VGND VPWR VPWR _08644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05856_ _05855_/Q _05887_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05173__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[12\].FF OVHB\[27\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[27\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08575_ _08574_/Q _08582_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05787_ _05799_/CLK line[11] VGND VGND VPWR VPWR _05788_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13390__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11903__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07526_ _07518_/CLK line[24] VGND VGND VPWR VPWR _07526_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08484__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _07457_/A _07462_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06408_ _06408_/CLK line[25] VGND VGND VPWR VPWR _06409_/A sky130_fd_sc_hd__dfxtp_1
X_07388_ _07380_/CLK line[89] VGND VGND VPWR VPWR _07388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09127_ _09127_/A _09142_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06339_ _06338_/Q _06342_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06732__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09058_ _09068_/CLK line[84] VGND VGND VPWR VPWR _09058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08009_ _08008_/Q _08022_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10254__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[9\].VALID\[3\].FF OVHB\[9\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[9\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05348__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11020_ _11002_/CLK line[85] VGND VGND VPWR VPWR _11020_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08302__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[14\].FF OVHB\[17\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[17\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13565__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08659__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07563__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08021__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12971_ _12970_/Q _12992_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11922_ _11934_/CLK line[113] VGND VGND VPWR VPWR _11923_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05083__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _11853_/A _11872_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11813__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[3\]_A0 _11402_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10804_ _10804_/CLK line[114] VGND VGND VPWR VPWR _10804_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06907__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11784_ _11776_/CLK line[50] VGND VGND VPWR VPWR _11785_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04920__B2 _04920_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05811__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13523_ _13522_/Q _13552_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10429__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10735_ _10734_/Q _10752_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[8\].VALID\[14\].TOBUF OVHB\[8\].VALID\[14\].FF/Q OVHB\[8\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_10666_ _10656_/CLK line[51] VGND VGND VPWR VPWR _10667_/A sky130_fd_sc_hd__dfxtp_1
X_13454_ _13468_/CLK line[60] VGND VGND VPWR VPWR _13454_/Q sky130_fd_sc_hd__dfxtp_1
X_12405_ _12405_/A _12432_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
X_13385_ _13384_/Q _13412_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_10597_ _10596_/Q _10612_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07738__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12336_ _12352_/CLK line[61] VGND VGND VPWR VPWR _12336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10164__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12267_ _12267_/A _12292_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05258__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11218_ _11216_/CLK line[62] VGND VGND VPWR VPWR _11218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12198_ _12204_/CLK line[126] VGND VGND VPWR VPWR _12199_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[21\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11149_ _11149_/A _11172_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07473__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[7\].VALID\[5\].FF OVHB\[7\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[7\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05710_ _05710_/CLK _05711_/X VGND VGND VPWR VPWR _05708_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[28\].VALID\[10\].TOBUF OVHB\[28\].VALID\[10\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06089__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06690_ _06690_/CLK _06691_/X VGND VGND VPWR VPWR _06682_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[1\].VALID\[13\].TOBUF OVHB\[1\].VALID\[13\].FF/Q OVHB\[1\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05571__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05641_ _13909_/X wr VGND VGND VPWR VPWR _05641_/X sky130_fd_sc_hd__and2_1
XFILLER_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08360_ _08358_/CLK line[21] VGND VGND VPWR VPWR _08361_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[9\].TOBUF OVHB\[10\].VALID\[9\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
X_05572_ _13909_/X VGND VGND VPWR VPWR _05572_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05721__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07311_ _07310_/Q _07322_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDATA\[6\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _12990_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10339__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08291_ _08290_/Q _08302_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07242_ _07232_/CLK line[22] VGND VGND VPWR VPWR _07242_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04915__A A_h[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07173_ _07172_/Q _07182_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12554__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07648__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06124_ _06108_/CLK line[23] VGND VGND VPWR VPWR _06125_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12851__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06055_ _06054_/Q _06062_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09863__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05746__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05006_ _05000_/CLK line[24] VGND VGND VPWR VPWR _05006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09814_ _09834_/CLK line[60] VGND VGND VPWR VPWR _09814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10802__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A _09772_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06957_ _06956_/Q _06972_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_05908_ _05902_/CLK line[52] VGND VGND VPWR VPWR _05909_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06888_ _06892_/CLK line[116] VGND VGND VPWR VPWR _06888_/Q sky130_fd_sc_hd__dfxtp_1
X_09676_ _09694_/CLK line[125] VGND VGND VPWR VPWR _09677_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05839_ _05838_/Q _05852_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_08627_ _08626_/Q _08652_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08560_/CLK line[126] VGND VGND VPWR VPWR _08559_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08792__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09103__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[7\].FF OVHB\[5\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[5\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ _07509_/A _07532_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_08489_ _08488_/Q _08512_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _10520_/CLK line[127] VGND VGND VPWR VPWR _10521_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10451_ _10451_/A _10472_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[5\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _12605_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06462__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13170_ _13194_/CLK line[58] VGND VGND VPWR VPWR _13170_/Q sky130_fd_sc_hd__dfxtp_1
X_10382_ _10384_/CLK line[49] VGND VGND VPWR VPWR _10382_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12121_ _12120_/Q _12152_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09773__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05078__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12052_ _12072_/CLK line[59] VGND VGND VPWR VPWR _12052_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13295__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11003_ _11002_/Q _11032_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[10\].FF OVHB\[23\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[23\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[4\].TOBUF OVHB\[19\].VALID\[4\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08389__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08967__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08686__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12954_ _12953_/Q _12957_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_11905_ _11905_/CLK _11906_/X VGND VGND VPWR VPWR _11901_/CLK sky130_fd_sc_hd__dlclkp_1
X_12885_ _12885_/CLK _12886_/X VGND VGND VPWR VPWR _12881_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11543__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06637__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11836_ _11872_/A wr VGND VGND VPWR VPWR _11836_/X sky130_fd_sc_hd__and2_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09013__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].CGAND_A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[25\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _09945_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11767_ _11872_/A VGND VGND VPWR VPWR _11767_/Y sky130_fd_sc_hd__inv_2
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09948__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13506_ _13506_/A _13517_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10718_ _10728_/CLK line[80] VGND VGND VPWR VPWR _10718_/Q sky130_fd_sc_hd__dfxtp_1
X_11698_ _11706_/CLK line[16] VGND VGND VPWR VPWR _11698_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07111__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13437_ _13439_/CLK line[38] VGND VGND VPWR VPWR _13437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[13\].VALID\[12\].FF OVHB\[13\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[13\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10649_ _10648_/Q _10682_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
X_13368_ _13368_/A _13377_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[9\].FF OVHB\[3\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[3\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12319_ _12311_/CLK line[39] VGND VGND VPWR VPWR _12320_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10472__A _13931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13299_ _13285_/CLK line[103] VGND VGND VPWR VPWR _13300_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10191__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11718__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07860_ _07854_/CLK line[63] VGND VGND VPWR VPWR _07860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06811_ _06811_/A _06832_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07791_ _07790_/Q _07812_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06742_ _06740_/CLK line[49] VGND VGND VPWR VPWR _06742_/Q sky130_fd_sc_hd__dfxtp_1
X_09530_ _09554_/CLK line[58] VGND VGND VPWR VPWR _09530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[0\].TOBUF OVHB\[0\].VALID\[0\].FF/Q OVHB\[0\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_09461_ _09460_/Q _09492_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06673_ _06673_/A _06692_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11453__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05624_ _05632_/CLK line[50] VGND VGND VPWR VPWR _05624_/Q sky130_fd_sc_hd__dfxtp_1
X_08412_ _08410_/CLK line[59] VGND VGND VPWR VPWR _08412_/Q sky130_fd_sc_hd__dfxtp_1
X_09392_ _09414_/CLK line[123] VGND VGND VPWR VPWR _09392_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[3\].TOBUF OVHB\[25\].VALID\[3\].FF/Q OVHB\[25\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__05451__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10069__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08343_ _08342_/Q _08372_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05555_ _05554_/Q _05572_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10647__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08274_ _08282_/CLK line[124] VGND VGND VPWR VPWR _08274_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08762__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05486_ _05476_/CLK line[115] VGND VGND VPWR VPWR _05487_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10366__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07225_ _07224_/Q _07252_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13958__A A_h[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12284__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[31\].VALID\[3\].FF OVHB\[31\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[31\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _09560_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07378__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07156_ _07170_/CLK line[125] VGND VGND VPWR VPWR _07156_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[30\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06107_ _06107_/A _06132_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07087_ _07086_/Q _07112_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09593__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06038_ _06050_/CLK line[126] VGND VGND VPWR VPWR _06038_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11628__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10532__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05626__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08002__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13843__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07989_ _07989_/A _08022_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08937__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09728_ _09727_/Q _09737_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07841__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12459__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09659_ _09659_/CLK line[103] VGND VGND VPWR VPWR _09660_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11941__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12669_/Q _12677_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11605_/CLK line[104] VGND VGND VPWR VPWR _11621_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[24\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[0\]_A3 _13554_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[9\].TOBUF OVHB\[17\].VALID\[9\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _11552_/A _11557_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _10473_/CLK line[105] VGND VGND VPWR VPWR _10504_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12194__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11483_ _11479_/CLK line[41] VGND VGND VPWR VPWR _11483_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10707__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07288__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06192__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13222_ _13221_/Q _13237_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
X_10434_ _10433_/Q _10437_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[2\].TOBUF OVHB\[31\].VALID\[2\].FF/Q OVHB\[31\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10365_ _10365_/CLK _10366_/X VGND VGND VPWR VPWR _10341_/CLK sky130_fd_sc_hd__dlclkp_1
X_13153_ _13163_/CLK line[36] VGND VGND VPWR VPWR _13153_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[14\].FF OVHB\[8\].V/CLK A[23] VGND VGND VPWR VPWR OVHB\[8\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[12\].VALID\[1\].FF OVHB\[12\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[12\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12104_ _12103_/Q _12117_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[23\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _09175_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_88_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13084_ _13083_/Q _13097_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_10296_ _13931_/X wr VGND VGND VPWR VPWR _10296_/X sky130_fd_sc_hd__and2_1
X_12035_ _12019_/CLK line[37] VGND VGND VPWR VPWR _12035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10442__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[13\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _06305_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[18\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12012__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13986_ _13982_/X _13990_/B _13990_/A _13990_/D VGND VGND VPWR VPWR _13986_/X sky130_fd_sc_hd__and4b_4
XANTENNA__07751__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12369__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12937_ _12937_/CLK line[65] VGND VGND VPWR VPWR _12937_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11273__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06367__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12868_ _12867_/Q _12887_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_11819_ _11823_/CLK line[66] VGND VGND VPWR VPWR _11820_/A sky130_fd_sc_hd__dfxtp_1
X_12799_ _12803_/CLK line[2] VGND VGND VPWR VPWR _12799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09678__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05340_ _05332_/CLK line[63] VGND VGND VPWR VPWR _05341_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10617__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05271_ _05270_/Q _05292_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07010_ _07030_/CLK line[58] VGND VGND VPWR VPWR _07010_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07776__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12832__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07926__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[6\].FF OVHB\[28\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[28\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08961_ _08947_/CLK line[40] VGND VGND VPWR VPWR _08961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[8\].TOBUF OVHB\[23\].VALID\[8\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11448__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07912_ _07912_/A _07917_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
X_08892_ _08891_/Q _08897_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07843_ _07837_/CLK line[41] VGND VGND VPWR VPWR _07843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[3\].FF OVHB\[10\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[10\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07774_ _07774_/A _07777_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
X_04986_ _05000_/CLK line[29] VGND VGND VPWR VPWR _04987_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[12\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _05920_/CLK sky130_fd_sc_hd__clkbuf_4
X_09513_ _09507_/CLK line[36] VGND VGND VPWR VPWR _09513_/Q sky130_fd_sc_hd__dfxtp_1
X_06725_ _06725_/CLK _06726_/X VGND VGND VPWR VPWR _06711_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_65_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11183__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06277__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06656_ _06832_/A wr VGND VGND VPWR VPWR _06656_/X sky130_fd_sc_hd__and2_1
X_09444_ _09443_/Q _09457_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05181__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05607_ _13909_/X VGND VGND VPWR VPWR _05607_/Y sky130_fd_sc_hd__inv_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09375_ _09365_/CLK line[101] VGND VGND VPWR VPWR _09375_/Q sky130_fd_sc_hd__dfxtp_1
X_06587_ _06551_/A VGND VGND VPWR VPWR _06587_/Y sky130_fd_sc_hd__inv_2
XANTENNA_MUX.MUX\[31\]_A2 _11851_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08326_ _08325_/Q _08337_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08492__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05538_ _05568_/CLK line[16] VGND VGND VPWR VPWR _05538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08257_ _08257_/CLK line[102] VGND VGND VPWR VPWR _08258_/A sky130_fd_sc_hd__dfxtp_1
X_05469_ _05468_/Q _05502_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07208_ _07208_/A _07217_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_08188_ _08187_/Q _08197_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07139_ _07117_/CLK line[103] VGND VGND VPWR VPWR _07139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06740__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10150_ _10149_/Q _10157_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11358__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10081_ _10073_/CLK line[40] VGND VGND VPWR VPWR _10082_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].CGAND _12151_/A wr VGND VGND VPWR VPWR OVHB\[3\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__05356__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[9\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13573__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13840_ _13839_/Q _13867_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08667__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[8\].FF OVHB\[26\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[26\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13771_ _13763_/CLK line[77] VGND VGND VPWR VPWR _13771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10983_ _10977_/CLK line[68] VGND VGND VPWR VPWR _10983_/Q sky130_fd_sc_hd__dfxtp_1
X_12722_ _12721_/Q _12747_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05091__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[0\].TOBUF OVHB\[7\].VALID\[0\].FF/Q OVHB\[7\].INV/Y VGND VGND VPWR
+ VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09141__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _12667_/CLK line[78] VGND VGND VPWR VPWR _12653_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _05535_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11604_ _11603_/Q _11627_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06915__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12583_/Q _12607_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _11535_/CLK line[79] VGND VGND VPWR VPWR _11535_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11466_ _11466_/A _11487_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[16\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13748__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13205_ _13213_/CLK line[74] VGND VGND VPWR VPWR _13205_/Q sky130_fd_sc_hd__dfxtp_1
X_10417_ _10405_/CLK line[65] VGND VGND VPWR VPWR _10418_/A sky130_fd_sc_hd__dfxtp_1
X_11397_ _11395_/CLK line[1] VGND VGND VPWR VPWR _11397_/Q sky130_fd_sc_hd__dfxtp_1
X_13136_ _13135_/Q _13167_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
X_10348_ _10347_/Q _10367_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10172__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13067_ _13075_/CLK line[11] VGND VGND VPWR VPWR _13067_/Q sky130_fd_sc_hd__dfxtp_1
X_10279_ _10277_/CLK line[2] VGND VGND VPWR VPWR _10279_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05266__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12018_ _12017_/Q _12047_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09316__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13483__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07481__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[13\].INV _13955_/X VGND VGND VPWR VPWR OVHB\[13\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12099__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13969_ A_h[4] VGND VGND VPWR VPWR _13979_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12677__A _12712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06510_ _06509_/Q _06517_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[13\].TOBUF OVHB\[14\].VALID\[13\].FF/Q OVHB\[14\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
X_07490_ _07489_/Q _07497_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12396__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06441_ _06421_/CLK line[40] VGND VGND VPWR VPWR _06441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[28\].INV _13976_/X VGND VGND VPWR VPWR OVHB\[28\].INV/Y sky130_fd_sc_hd__inv_2
X_09160_ _09159_/Q _09177_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_06372_ _06371_/Q _06377_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[12\].FF OVHB\[4\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[4\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08111_ _08113_/CLK line[35] VGND VGND VPWR VPWR _08112_/A sky130_fd_sc_hd__dfxtp_1
X_05323_ _05299_/CLK line[41] VGND VGND VPWR VPWR _05324_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10347__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09091_ _09085_/CLK line[99] VGND VGND VPWR VPWR _09091_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08042_ _08041_/Q _08057_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_05254_ _05253_/Q _05257_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13658__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12562__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05185_ _05185_/CLK _05186_/X VGND VGND VPWR VPWR _05157_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07656__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09993_ _10011_/CLK line[14] VGND VGND VPWR VPWR _09993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ _08943_/Q _08967_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09871__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08875_ _08869_/CLK line[15] VGND VGND VPWR VPWR _08875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13971__A A_h[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10810__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07826_ _07825_/Q _07847_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05904__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07757_ _07773_/CLK line[1] VGND VGND VPWR VPWR _07757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04969_ _04947_/CLK line[7] VGND VGND VPWR VPWR _04969_/Q sky130_fd_sc_hd__dfxtp_1
X_06708_ _06708_/A _06727_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_07688_ _07687_/Q _07707_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12737__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[31\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09427_ _09427_/CLK line[11] VGND VGND VPWR VPWR _09428_/A sky130_fd_sc_hd__dfxtp_1
X_06639_ _06633_/CLK line[2] VGND VGND VPWR VPWR _06639_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].INV_A _13972_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09358_ _09357_/Q _09387_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XMUX.MUX\[12\] _10830_/Z _05020_/Z _13490_/Z _06840_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[12] sky130_fd_sc_hd__mux4_1
X_08309_ _08329_/CLK line[12] VGND VGND VPWR VPWR _08309_/Q sky130_fd_sc_hd__dfxtp_1
X_09289_ _09307_/CLK line[76] VGND VGND VPWR VPWR _09289_/Q sky130_fd_sc_hd__dfxtp_1
X_11320_ _11319_/Q _11347_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[28\].VALID\[10\].FF OVHB\[28\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[28\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12472__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11251_ _11251_/CLK line[77] VGND VGND VPWR VPWR _11251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ _10201_/Q _10227_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06470__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11182_ _11181_/Q _11207_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11088__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10133_ _10145_/CLK line[78] VGND VGND VPWR VPWR _10134_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[5\].TOBUF OVHB\[5\].VALID\[5\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09781__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10064_ _10063_/Q _10087_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08397__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10720__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13823_ _13822_/Q _13832_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13754_ _13746_/CLK line[55] VGND VGND VPWR VPWR _13754_/Q sky130_fd_sc_hd__dfxtp_1
X_10966_ _10965_/Q _10997_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[12\].FF OVHB\[18\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[18\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12705_ _12704_/Q _12712_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12647__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11551__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13685_ _13684_/Q _13692_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_10897_ _10903_/CLK line[43] VGND VGND VPWR VPWR _10897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _12638_/CLK line[56] VGND VGND VPWR VPWR _12636_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06645__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12567_ _12566_/Q _12572_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09956__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11518_ _11500_/CLK line[57] VGND VGND VPWR VPWR _11518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12498_ _12490_/CLK line[121] VGND VGND VPWR VPWR _12498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13478__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11449_ _11449_/A _11452_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06380__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13119_ _13118_/Q _13132_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
X_06990_ _06990_/A _07007_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[21\]_A1 _10391_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05941_ _05929_/CLK line[67] VGND VGND VPWR VPWR _05941_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11726__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08660_ _08659_/Q _08687_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_05872_ _05872_/A _05887_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07611_ _07633_/CLK line[77] VGND VGND VPWR VPWR _07611_/Q sky130_fd_sc_hd__dfxtp_1
X_08591_ _08609_/CLK line[13] VGND VGND VPWR VPWR _08591_/Q sky130_fd_sc_hd__dfxtp_1
X_07542_ _07541_/Q _07567_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[0\].TOBUF OVHB\[12\].VALID\[0\].FF/Q OVHB\[12\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
X_07473_ _07467_/CLK line[14] VGND VGND VPWR VPWR _07473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11461__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09212_ _09352_/A VGND VGND VPWR VPWR _09212_/Y sky130_fd_sc_hd__inv_2
X_06424_ _06423_/Q _06447_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06555__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10077__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06355_ _06353_/CLK line[15] VGND VGND VPWR VPWR _06356_/A sky130_fd_sc_hd__dfxtp_1
X_09143_ _09147_/CLK line[0] VGND VGND VPWR VPWR _09143_/Q sky130_fd_sc_hd__dfxtp_1
X_05306_ _05305_/Q _05327_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_09074_ _09073_/Q _09107_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08770__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06286_ _06286_/A _06307_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13388__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08025_ _08033_/CLK line[10] VGND VGND VPWR VPWR _08025_/Q sky130_fd_sc_hd__dfxtp_1
X_05237_ _05253_/CLK line[1] VGND VGND VPWR VPWR _05238_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07386__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05168_ _05168_/A _05187_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[10\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11486__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09976_ _09978_/CLK line[120] VGND VGND VPWR VPWR _09977_/A sky130_fd_sc_hd__dfxtp_1
X_05099_ _05093_/CLK line[66] VGND VGND VPWR VPWR _05099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08927_ _08926_/Q _08932_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11636__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[3\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _12220_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_131_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08858_ _08850_/CLK line[121] VGND VGND VPWR VPWR _08859_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05634__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[10\].FF OVHB\[0\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[0\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08010__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07809_ _07808_/Q _07812_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08789_ _08789_/A _08792_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13851__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10820_ _10820_/CLK _10821_/X VGND VGND VPWR VPWR _10804_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_77_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08945__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10751_ _13932_/X wr VGND VGND VPWR VPWR _10751_/X sky130_fd_sc_hd__and2_1
XANTENNA_DATA\[3\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13470_ _13468_/CLK line[53] VGND VGND VPWR VPWR _13470_/Q sky130_fd_sc_hd__dfxtp_1
X_10682_ _13932_/X VGND VGND VPWR VPWR _10682_/Y sky130_fd_sc_hd__inv_2
X_12421_ _12420_/Q _12432_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_12352_ _12352_/CLK line[54] VGND VGND VPWR VPWR _12352_/Q sky130_fd_sc_hd__dfxtp_1
X_11303_ _11303_/A _11312_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
X_12283_ _12282_/Q _12292_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07296__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05809__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11234_ _11216_/CLK line[55] VGND VGND VPWR VPWR _11235_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11165_ _11164_/Q _11172_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10116_ _10100_/CLK line[56] VGND VGND VPWR VPWR _10116_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[10\].TOBUF OVHB\[8\].VALID\[10\].FF/Q OVHB\[8\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_11096_ _11090_/CLK line[120] VGND VGND VPWR VPWR _11096_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10450__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10047_ _10047_/A _10052_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].CG clk OVHB\[16\].CGAND/X VGND VGND VPWR VPWR OVHB\[16\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05544__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13806_ _13822_/CLK line[93] VGND VGND VPWR VPWR _13806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[2\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _11275_/CLK sky130_fd_sc_hd__clkbuf_4
X_11998_ _12002_/CLK line[20] VGND VGND VPWR VPWR _11998_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _13736_/Q _13762_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12377__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10949_ _10948_/Q _10962_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
X_13668_ _13682_/CLK line[30] VGND VGND VPWR VPWR _13669_/A sky130_fd_sc_hd__dfxtp_1
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12619_ _12618_/Q _12642_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
X_13599_ _13598_/Q _13622_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09686__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06140_ _06140_/A _06167_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10625__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06071_ _06077_/CLK line[13] VGND VGND VPWR VPWR _06071_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13001__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05719__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05022_ _05022_/A _05047_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[5\].TOBUF OVHB\[10\].VALID\[5\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XDEC.DEC0.AND2 A[7] A[8] VGND VGND VPWR VPWR _13923_/D sky130_fd_sc_hd__and2b_2
X_09830_ _09834_/CLK line[53] VGND VGND VPWR VPWR _09830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12840__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07934__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09761_ _09760_/Q _09772_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_06973_ _07001_/CLK line[32] VGND VGND VPWR VPWR _06973_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[10\].FF OVHB\[14\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[14\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08712_ _08710_/CLK line[54] VGND VGND VPWR VPWR _08712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[29\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05924_ _05923_/Q _05957_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_09692_ _09694_/CLK line[118] VGND VGND VPWR VPWR _09692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08643_ _08643_/A _08652_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05855_ _05871_/CLK line[42] VGND VGND VPWR VPWR _05855_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13026__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _08560_/CLK line[119] VGND VGND VPWR VPWR _08574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05786_ _05785_/Q _05817_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _07524_/Q _07532_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06285__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07456_ _07446_/CLK line[120] VGND VGND VPWR VPWR _07457_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[1\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _08090_/CLK sky130_fd_sc_hd__clkbuf_4
X_06407_ _06406_/Q _06412_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
X_07387_ _07387_/A _07392_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09126_ _09116_/CLK line[115] VGND VGND VPWR VPWR _09127_/A sky130_fd_sc_hd__dfxtp_1
X_06338_ _06320_/CLK line[121] VGND VGND VPWR VPWR _06338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04932__A2_N _04932_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _09057_/A _09072_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06269_ _06268_/Q _06272_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_08008_ _08000_/CLK line[116] VGND VGND VPWR VPWR _08008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12750__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ _09958_/Q _09982_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11366__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _12962_/CLK line[95] VGND VGND VPWR VPWR _12970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11921_ _11920_/Q _11942_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13581__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11852_ _11846_/CLK line[81] VGND VGND VPWR VPWR _11853_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08675__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[21\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _08790_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_MUX.MUX\[3\]_A1 _05592_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10803_ _10802_/Q _10822_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_11783_ _11782_/Q _11802_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13522_ _13528_/CLK line[91] VGND VGND VPWR VPWR _13522_/Q sky130_fd_sc_hd__dfxtp_1
X_10734_ _10728_/CLK line[82] VGND VGND VPWR VPWR _10734_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[0\].TOBUF OVHB\[19\].VALID\[0\].FF/Q OVHB\[19\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DECH.DEC0.AND0_A A_h[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[11\]_A0 _04948_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13453_ _13453_/A _13482_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12925__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10665_ _10664_/Q _10682_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12404_ _12414_/CLK line[92] VGND VGND VPWR VPWR _12405_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06923__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13384_ _13394_/CLK line[28] VGND VGND VPWR VPWR _13384_/Q sky130_fd_sc_hd__dfxtp_1
X_10596_ _10594_/CLK line[19] VGND VGND VPWR VPWR _10596_/Q sky130_fd_sc_hd__dfxtp_1
X_12335_ _12334_/Q _12362_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[1\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12266_ _12268_/CLK line[29] VGND VGND VPWR VPWR _12267_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13756__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[11\].TOBUF OVHB\[24\].VALID\[11\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_11217_ _11216_/Q _11242_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
X_12197_ _12196_/Q _12222_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
X_11148_ _11148_/CLK line[30] VGND VGND VPWR VPWR _11149_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10180__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05274__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11079_ _11078_/Q _11102_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05852__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13491__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[12\].FF OVHB\[9\].V/CLK A[21] VGND VGND VPWR VPWR OVHB\[9\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05571__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05640_ _05640_/CLK _05641_/X VGND VGND VPWR VPWR _05632_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08585__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05571_ _13909_/X wr VGND VGND VPWR VPWR _05571_/X sky130_fd_sc_hd__and2_1
X_07310_ _07292_/CLK line[53] VGND VGND VPWR VPWR _07310_/Q sky130_fd_sc_hd__dfxtp_1
X_08290_ _08282_/CLK line[117] VGND VGND VPWR VPWR _08290_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[20\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _08405_/CLK sky130_fd_sc_hd__clkbuf_4
X_07241_ _07240_/Q _07252_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06833__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07172_ _07170_/CLK line[118] VGND VGND VPWR VPWR _07172_/Q sky130_fd_sc_hd__dfxtp_1
X_06123_ _06123_/A _06132_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10355__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05449__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06054_ _06050_/CLK line[119] VGND VGND VPWR VPWR _06054_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13666__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05005_ _05005_/A _05012_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05746__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07664__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09813_ _09812_/Q _09842_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10090__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09744_ _09760_/CLK line[28] VGND VGND VPWR VPWR _09745_/A sky130_fd_sc_hd__dfxtp_1
X_06956_ _06960_/CLK line[19] VGND VGND VPWR VPWR _06956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05907_ _05906_/Q _05922_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09675_ _09674_/Q _09702_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_06887_ _06886_/Q _06902_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11914__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08626_ _08646_/CLK line[29] VGND VGND VPWR VPWR _08626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05838_ _05836_/CLK line[20] VGND VGND VPWR VPWR _05838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05912__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08556_/Q _08582_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05769_ _05769_/A _05782_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07508_ _07518_/CLK line[30] VGND VGND VPWR VPWR _07509_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08488_ _08480_/CLK line[94] VGND VGND VPWR VPWR _08488_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07439_ _07438_/Q _07462_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[4\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07839__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[1\].FF OVHB\[20\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[20\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10450_ _10466_/CLK line[95] VGND VGND VPWR VPWR _10451_/A sky130_fd_sc_hd__dfxtp_1
X_09109_ _09109_/A _09142_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10265__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10381_ _10380_/Q _10402_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _12130_/CLK line[90] VGND VGND VPWR VPWR _12120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12480__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _12050_/Q _12082_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07574__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11002_ _11002_/CLK line[91] VGND VGND VPWR VPWR _11002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11096__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[5\].TOBUF OVHB\[17\].VALID\[5\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ _12937_/CLK line[73] VGND VGND VPWR VPWR _12953_/Q sky130_fd_sc_hd__dfxtp_1
X_11904_ _11903_/Q _11907_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
X_12884_ _12883_/Q _12887_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05822__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11835_ _11835_/CLK _11836_/X VGND VGND VPWR VPWR _11823_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_14_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[3\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[22\].CGAND_A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11766_ _11872_/A wr VGND VGND VPWR VPWR _11766_/X sky130_fd_sc_hd__and2_1
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13505_ _13497_/CLK line[69] VGND VGND VPWR VPWR _13506_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[2\].FF OVHB\[19\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[19\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _13932_/X VGND VGND VPWR VPWR _10717_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12655__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11872_/A VGND VGND VPWR VPWR _11697_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07749__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].CGAND_A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07111__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13436_ _13436_/A _13447_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06653__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10648_ _10656_/CLK line[48] VGND VGND VPWR VPWR _10648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ _13347_/CLK line[6] VGND VGND VPWR VPWR _13368_/A sky130_fd_sc_hd__dfxtp_1
X_10579_ _10579_/A _10612_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09964__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12318_ _12317_/Q _12327_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13298_ _13297_/Q _13307_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10903__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12249_ _12227_/CLK line[7] VGND VGND VPWR VPWR _12249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06810_ _06802_/CLK line[95] VGND VGND VPWR VPWR _06811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07790_ _07788_/CLK line[31] VGND VGND VPWR VPWR _07790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06741_ _06740_/Q _06762_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06828__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09460_ _09482_/CLK line[26] VGND VGND VPWR VPWR _09460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06672_ _06682_/CLK line[17] VGND VGND VPWR VPWR _06673_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09204__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08411_ _08411_/A _08442_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
X_05623_ _05623_/A _05642_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
X_09391_ _09390_/Q _09422_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[4\].TOBUF OVHB\[23\].VALID\[4\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
X_08342_ _08358_/CLK line[27] VGND VGND VPWR VPWR _08342_/Q sky130_fd_sc_hd__dfxtp_1
X_05554_ _05568_/CLK line[18] VGND VGND VPWR VPWR _05554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05485_ _05484_/Q _05502_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_08273_ _08272_/Q _08302_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06563__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07224_ _07232_/CLK line[28] VGND VGND VPWR VPWR _07224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07155_ _07155_/A _07182_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05179__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06106_ _06108_/CLK line[29] VGND VGND VPWR VPWR _06107_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07086_ _07098_/CLK line[93] VGND VGND VPWR VPWR _07086_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[4\].FF OVHB\[17\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[17\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13396__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06037_ _06036_/Q _06062_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[5\].VALID\[10\].FF OVHB\[5\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[5\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07988_ _08000_/CLK line[112] VGND VGND VPWR VPWR _07989_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ _09721_/CLK line[6] VGND VGND VPWR VPWR _09727_/Q sky130_fd_sc_hd__dfxtp_1
X_06939_ _06938_/Q _06972_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11644__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06738__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09658_ _09657_/Q _09667_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09114__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08609_ _08609_/CLK line[7] VGND VGND VPWR VPWR _08610_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11941__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09577_/CLK line[71] VGND VGND VPWR VPWR _09590_/A sky130_fd_sc_hd__dfxtp_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11619_/Q _11627_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _11535_/CLK line[72] VGND VGND VPWR VPWR _11552_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ _10501_/Q _10507_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11482_ _11482_/A _11487_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _13213_/CLK line[67] VGND VGND VPWR VPWR _13221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10433_ _10405_/CLK line[73] VGND VGND VPWR VPWR _10433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05089__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13152_ _13152_/A _13167_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
X_10364_ _10363_/Q _10367_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11819__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12103_ _12109_/CLK line[68] VGND VGND VPWR VPWR _12103_/Q sky130_fd_sc_hd__dfxtp_1
X_13083_ _13075_/CLK line[4] VGND VGND VPWR VPWR _13083_/Q sky130_fd_sc_hd__dfxtp_1
X_10295_ _10295_/CLK _10296_/X VGND VGND VPWR VPWR _10277_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07882__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12034_ _12033_/Q _12047_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[6\].FF OVHB\[15\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[15\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13985_ _13982_/X _13990_/A _13990_/B _13990_/D VGND VGND VPWR VPWR _13985_/X sky130_fd_sc_hd__and4bb_4
XANTENNA_DATA\[24\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12936_ _12935_/Q _12957_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05552__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12867_ _12881_/CLK line[33] VGND VGND VPWR VPWR _12867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08863__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11818_ _11817_/Q _11837_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ _12797_/Q _12817_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12385__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11749_ _11757_/CLK line[34] VGND VGND VPWR VPWR _11750_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07479__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05270_ _05278_/CLK line[31] VGND VGND VPWR VPWR _05270_/Q sky130_fd_sc_hd__dfxtp_1
X_13419_ _13439_/CLK line[44] VGND VGND VPWR VPWR _13419_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07776__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09694__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[10\].FF OVHB\[19\].V/CLK A[19] VGND VGND VPWR VPWR OVHB\[19\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10633__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08960_ _08960_/A _08967_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05727__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07911_ _07905_/CLK line[72] VGND VGND VPWR VPWR _07912_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[9\].TOBUF OVHB\[21\].VALID\[9\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08103__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08891_ _08869_/CLK line[8] VGND VGND VPWR VPWR _08891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07842_ _07842_/A _07847_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07942__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06201__A _06272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07773_ _07773_/CLK line[9] VGND VGND VPWR VPWR _07774_/A sky130_fd_sc_hd__dfxtp_1
X_04985_ _04984_/Q _05012_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_09512_ _09511_/Q _09527_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06724_ _06723_/Q _06727_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09443_ _09427_/CLK line[4] VGND VGND VPWR VPWR _09443_/Q sky130_fd_sc_hd__dfxtp_1
X_06655_ _06655_/CLK _06656_/X VGND VGND VPWR VPWR _06633_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09869__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05606_ _13909_/X wr VGND VGND VPWR VPWR _05606_/X sky130_fd_sc_hd__and2_1
X_09374_ _09373_/Q _09387_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[13\].VALID\[8\].FF OVHB\[13\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[13\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06586_ _06551_/A wr VGND VGND VPWR VPWR _06586_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.MUX\[31\]_A3 _13601_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12295__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08325_ _08329_/CLK line[5] VGND VGND VPWR VPWR _08325_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13969__A A_h[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10808__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05537_ _13909_/X VGND VGND VPWR VPWR _05537_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06293__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08256_ _08255_/Q _08267_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
X_05468_ _05476_/CLK line[112] VGND VGND VPWR VPWR _05468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07207_ _07183_/CLK line[6] VGND VGND VPWR VPWR _07208_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08187_ _08175_/CLK line[70] VGND VGND VPWR VPWR _08187_/Q sky130_fd_sc_hd__dfxtp_1
X_05399_ _05398_/Q _05432_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
X_07138_ _07137_/Q _07147_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10543__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07069_ _07043_/CLK line[71] VGND VGND VPWR VPWR _07069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10080_ _10080_/A _10087_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07852__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11374__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06468__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13770_ _13769_/Q _13797_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10982_ _10982_/A _10997_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12721_ _12741_/CLK line[109] VGND VGND VPWR VPWR _12721_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09422__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09779__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09141__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12652_ _12652_/A _12677_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[1\].TOBUF OVHB\[5\].VALID\[1\].FF/Q OVHB\[5\].INV/Y VGND VGND VPWR
+ VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11603_ _11605_/CLK line[110] VGND VGND VPWR VPWR _11603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10718__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12583_ _12601_/CLK line[46] VGND VGND VPWR VPWR _12583_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _11534_/A _11557_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12933__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11465_ _11479_/CLK line[47] VGND VGND VPWR VPWR _11466_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05397__A _13908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _13203_/Q _13237_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_10416_ _10415_/Q _10437_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06931__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11396_ _11395_/Q _11417_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11549__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13135_ _13163_/CLK line[42] VGND VGND VPWR VPWR _13135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10347_ _10341_/CLK line[33] VGND VGND VPWR VPWR _10347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[11\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09019__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13066_ _13066_/A _13097_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_10278_ _10277_/Q _10297_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_12017_ _12019_/CLK line[43] VGND VGND VPWR VPWR _12017_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08858__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[14\].TOBUF OVHB\[10\].VALID\[14\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XANTENNA__09316__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11284__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06378__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13968_ _13958_/X _13964_/B _13960_/X _13966_/D VGND VGND VPWR VPWR _13968_/X sky130_fd_sc_hd__and4_4
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05282__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12919_ _12918_/Q _12922_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_13899_ _13898_/Q _13902_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[30\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _11660_/CLK sky130_fd_sc_hd__clkbuf_4
X_06440_ _06440_/A _06447_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08593__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[2\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06371_ _06353_/CLK line[8] VGND VGND VPWR VPWR _06371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08110_ _08109_/Q _08127_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_05322_ _05321_/Q _05327_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_09090_ _09089_/Q _09107_/Y VGND VGND VPWR VPWR _13570_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06691__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08041_ _08033_/CLK line[3] VGND VGND VPWR VPWR _08041_/Q sky130_fd_sc_hd__dfxtp_1
X_05253_ _05253_/CLK line[9] VGND VGND VPWR VPWR _05253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__04923__B _04923_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11102__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06841__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05184_ _05183_/Q _05187_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11459__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10363__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09992_ _09992_/A _10017_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05457__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08943_ _08947_/CLK line[46] VGND VGND VPWR VPWR _08943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[23\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13674__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08874_ _08873_/Q _08897_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08768__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07825_ _07837_/CLK line[47] VGND VGND VPWR VPWR _07825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07756_ _07756_/A _07777_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06866__A _06832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04968_ _04967_/Q _04977_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05192__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06707_ _06711_/CLK line[33] VGND VGND VPWR VPWR _06708_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07687_ _07679_/CLK line[97] VGND VGND VPWR VPWR _07687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11922__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09426_ _09426_/A _09457_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
X_06638_ _06637_/Q _06657_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[13\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09357_ _09365_/CLK line[107] VGND VGND VPWR VPWR _09357_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10538__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[1\].FF OVHB\[6\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[6\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06569_ _06565_/CLK line[98] VGND VGND VPWR VPWR _06570_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08308_ _08307_/Q _08337_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08008__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _09288_/A _09317_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13849__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08239_ _08257_/CLK line[108] VGND VGND VPWR VPWR _08239_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[14\].TOBUF OVHB\[30\].VALID\[14\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
X_11250_ _11250_/A _11277_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10201_ _10217_/CLK line[109] VGND VGND VPWR VPWR _10201_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10273__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11181_ _11191_/CLK line[45] VGND VGND VPWR VPWR _11181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__05367__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10132_ _10131_/Q _10157_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[6\].TOBUF OVHB\[3\].VALID\[6\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10063_ _10073_/CLK line[46] VGND VGND VPWR VPWR _10063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07582__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[9\].TOBUF OVHB\[28\].VALID\[9\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_21_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06198__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13822_ _13822_/CLK line[86] VGND VGND VPWR VPWR _13822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13753_ _13752_/Q _13762_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10965_ _10977_/CLK line[74] VGND VGND VPWR VPWR _10965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ _12708_/CLK line[87] VGND VGND VPWR VPWR _12704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13684_ _13682_/CLK line[23] VGND VGND VPWR VPWR _13684_/Q sky130_fd_sc_hd__dfxtp_1
X_10896_ _10895_/Q _10927_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05830__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _12634_/Q _12642_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10448__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[17\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12566_ _12560_/CLK line[24] VGND VGND VPWR VPWR _12566_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _11516_/Q _11522_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12663__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12497_ _12496_/Q _12502_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07757__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11448_ _11440_/CLK line[25] VGND VGND VPWR VPWR _11449_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[3\].FF OVHB\[4\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[4\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ _11378_/Q _11382_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09972__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13118_ _13120_/CLK line[20] VGND VGND VPWR VPWR _13118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08231__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_MUX.MUX\[21\]_A2 _13541_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10911__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05940_ _05939_/Q _05957_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_13049_ _13048_/Q _13062_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05871_ _05871_/CLK line[35] VGND VGND VPWR VPWR _05872_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07610_ _07610_/A _07637_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11592__A _11592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08590_ _08589_/Q _08617_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07541_ _07539_/CLK line[45] VGND VGND VPWR VPWR _07541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12838__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[1\].TOBUF OVHB\[10\].VALID\[1\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_07472_ _07471_/Q _07497_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09211_ _09352_/A wr VGND VGND VPWR VPWR _09211_/X sky130_fd_sc_hd__and2_1
X_06423_ _06421_/CLK line[46] VGND VGND VPWR VPWR _06423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[8\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09142_ _13923_/X VGND VGND VPWR VPWR _09142_/Y sky130_fd_sc_hd__inv_2
X_06354_ _06354_/A _06377_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08406__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].V_RESET_B rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05305_ _05299_/CLK line[47] VGND VGND VPWR VPWR _05305_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12573__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09073_ _09085_/CLK line[96] VGND VGND VPWR VPWR _09073_/Q sky130_fd_sc_hd__dfxtp_1
X_06285_ _06285_/CLK line[111] VGND VGND VPWR VPWR _06286_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06571__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08024_ _08023_/Q _08057_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_05236_ _05236_/A _05257_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11189__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11767__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05167_ _05157_/CLK line[97] VGND VGND VPWR VPWR _05168_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09882__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11486__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09975_ _09974_/Q _09982_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
X_05098_ _05097_/Q _05117_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13982__A A_h[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08926_ _08922_/CLK line[24] VGND VGND VPWR VPWR _08926_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08498__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[18\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[2\].VALID\[5\].FF OVHB\[2\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[2\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08857_ _08857_/A _08862_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07808_ _07788_/CLK line[25] VGND VGND VPWR VPWR _07808_/Q sky130_fd_sc_hd__dfxtp_1
X_08788_ _08762_/CLK line[89] VGND VGND VPWR VPWR _08789_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07739_ _07739_/A _07742_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12748__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__04932__B1 A_h[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11652__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06746__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10750_ _10750_/CLK _10751_/X VGND VGND VPWR VPWR _10728_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09122__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09409_ _09409_/A _09422_/Y VGND VGND VPWR VPWR _07169_/Z sky130_fd_sc_hd__ebufn_2
X_10681_ _13932_/X wr VGND VGND VPWR VPWR _10681_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[28\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12420_ _12414_/CLK line[85] VGND VGND VPWR VPWR _12420_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08961__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13579__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12351_ _12350_/Q _12362_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_11302_ _11302_/CLK line[86] VGND VGND VPWR VPWR _11303_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].INV _13954_/X VGND VGND VPWR VPWR OVHB\[12\].INV/Y sky130_fd_sc_hd__inv_2
X_12282_ _12268_/CLK line[22] VGND VGND VPWR VPWR _12282_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[11\].TOBUF OVHB\[4\].VALID\[11\].FF/Q OVHB\[4\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_11233_ _11232_/Q _11242_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05097__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11164_ _11148_/CLK line[23] VGND VGND VPWR VPWR _11164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11827__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10115_ _10114_/Q _10122_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[27\].INV _13975_/X VGND VGND VPWR VPWR OVHB\[27\].INV/Y sky130_fd_sc_hd__inv_2
X_11095_ _11094_/Q _11102_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10046_ _10042_/CLK line[24] VGND VGND VPWR VPWR _10047_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13805_ _13805_/A _13832_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11997_ _11996_/Q _12012_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11562__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13736_ _13746_/CLK line[61] VGND VGND VPWR VPWR _13736_/Q sky130_fd_sc_hd__dfxtp_1
X_10948_ _10930_/CLK line[52] VGND VGND VPWR VPWR _10948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05560__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[7\].FF OVHB\[0\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[0\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10178__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13667_ _13666_/Q _13692_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
X_10879_ _10878_/Q _10892_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13132__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12618_ _12638_/CLK line[62] VGND VGND VPWR VPWR _12618_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13598_ _13598_/CLK line[126] VGND VGND VPWR VPWR _13598_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13489__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12393__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12549_ _12548_/Q _12572_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07487__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06070_ _06069_/Q _06097_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05021_ _05041_/CLK line[45] VGND VGND VPWR VPWR _05022_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC.DEC0.AND3 A[8] A[7] VGND VGND VPWR VPWR _13934_/D sky130_fd_sc_hd__and2_2
XOVHB\[29\].VALID\[0\].FF OVHB\[29\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[29\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11737__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10641__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09760_ _09760_/CLK line[21] VGND VGND VPWR VPWR _09760_/Q sky130_fd_sc_hd__dfxtp_1
X_06972_ _07111_/A VGND VGND VPWR VPWR _06972_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08896__A _13923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05735__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08711_ _08711_/A _08722_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08111__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05923_ _05929_/CLK line[64] VGND VGND VPWR VPWR _05923_/Q sky130_fd_sc_hd__dfxtp_1
X_09691_ _09691_/A _09702_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[29\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13307__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08642_ _08646_/CLK line[22] VGND VGND VPWR VPWR _08643_/A sky130_fd_sc_hd__dfxtp_1
X_05854_ _05853_/Q _05887_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13026__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08573_ _08572_/Q _08582_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12568__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05785_ _05799_/CLK line[10] VGND VGND VPWR VPWR _05785_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07524_ _07518_/CLK line[23] VGND VGND VPWR VPWR _07524_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05470__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[8\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10088__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07455_ _07455_/A _07462_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06406_ _06408_/CLK line[24] VGND VGND VPWR VPWR _06406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07386_ _07380_/CLK line[88] VGND VGND VPWR VPWR _07387_/A sky130_fd_sc_hd__dfxtp_1
X_09125_ _09124_/Q _09142_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10816__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06337_ _06336_/Q _06342_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07397__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09056_ _09068_/CLK line[83] VGND VGND VPWR VPWR _09057_/A sky130_fd_sc_hd__dfxtp_1
X_06268_ _06244_/CLK line[89] VGND VGND VPWR VPWR _06268_/Q sky130_fd_sc_hd__dfxtp_1
X_08007_ _08007_/A _08022_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_05219_ _05218_/Q _05222_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_06199_ _06198_/Q _06202_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[13\].TOBUF OVHB\[27\].VALID\[13\].FF/Q OVHB\[27\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10551__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09958_ _09978_/CLK line[126] VGND VGND VPWR VPWR _09958_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05645__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08909_ _08908_/Q _08932_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
X_09889_ _09888_/Q _09912_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_11920_ _11934_/CLK line[127] VGND VGND VPWR VPWR _11920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07860__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[27\].VALID\[2\].FF OVHB\[27\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[27\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11851_ _11850_/Q _11872_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12478__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10802_ _10804_/CLK line[113] VGND VGND VPWR VPWR _10802_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06476__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[3\]_A2 _13502_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11782_ _11776_/CLK line[49] VGND VGND VPWR VPWR _11782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13521_ _13520_/Q _13552_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_10733_ _10732_/Q _10752_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10576__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09787__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DECH.DEC0.AND0_B A_h[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13452_ _13468_/CLK line[59] VGND VGND VPWR VPWR _13453_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[1\].TOBUF OVHB\[17\].VALID\[1\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_10664_ _10656_/CLK line[50] VGND VGND VPWR VPWR _10664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[11\]_A1 _05578_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12402_/Q _12432_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10726__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[12\].TOBUF OVHB\[20\].VALID\[12\].FF/Q OVHB\[20\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_13383_ _13383_/A _13412_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_10595_ _10595_/A _10612_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13102__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _12352_/CLK line[60] VGND VGND VPWR VPWR _12334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07100__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12941__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12265_ _12264_/Q _12292_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11216_ _11216_/CLK line[61] VGND VGND VPWR VPWR _11216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12196_ _12204_/CLK line[125] VGND VGND VPWR VPWR _12196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11147_ _11146_/Q _11172_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09027__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11078_ _11090_/CLK line[126] VGND VGND VPWR VPWR _11078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10029_ _10029_/A _10052_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11292__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06386__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05570_ _05570_/CLK _05571_/X VGND VGND VPWR VPWR _05568_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_44_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13719_ _13701_/CLK line[39] VGND VGND VPWR VPWR _13719_/Q sky130_fd_sc_hd__dfxtp_1
X_07240_ _07232_/CLK line[21] VGND VGND VPWR VPWR _07240_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[1\].FF_D A[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[4\].FF OVHB\[25\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[25\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13797__A _13907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07171_ _07170_/Q _07182_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06122_ _06108_/CLK line[22] VGND VGND VPWR VPWR _06123_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07010__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[19\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _07775_/CLK sky130_fd_sc_hd__clkbuf_4
X_06053_ _06052_/Q _06062_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05004_ _05000_/CLK line[23] VGND VGND VPWR VPWR _05005_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[23\].VALID\[0\].TOBUF OVHB\[23\].VALID\[0\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04940_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_28_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11467__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09812_ _09834_/CLK line[59] VGND VGND VPWR VPWR _09812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09743_ _09742_/Q _09772_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_06955_ _06955_/A _06972_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13682__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05906_ _05902_/CLK line[51] VGND VGND VPWR VPWR _05906_/Q sky130_fd_sc_hd__dfxtp_1
X_09674_ _09694_/CLK line[124] VGND VGND VPWR VPWR _09674_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08776__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06886_ _06892_/CLK line[115] VGND VGND VPWR VPWR _06886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08625_ _08624_/Q _08652_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_05837_ _05836_/Q _05852_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08560_/CLK line[125] VGND VGND VPWR VPWR _08556_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ _05756_/CLK line[116] VGND VGND VPWR VPWR _05769_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07507_ _07507_/A _07532_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08487_ _08487_/A _08512_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11930__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05699_ _05698_/Q _05712_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ _07446_/CLK line[126] VGND VGND VPWR VPWR _07438_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09400__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07369_ _07369_/A _07392_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09108_ _09116_/CLK line[112] VGND VGND VPWR VPWR _09109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08016__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10380_ _10384_/CLK line[63] VGND VGND VPWR VPWR _10380_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13857__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09039_ _09038_/Q _09072_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12116__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[6\].FF OVHB\[23\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[23\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12050_ _12072_/CLK line[58] VGND VGND VPWR VPWR _12050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11001_ _11000_/Q _11032_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10281__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05375__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[15\].VALID\[6\].TOBUF OVHB\[15\].VALID\[6\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__13592__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12952_ _12951_/Q _12957_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07590__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11903_ _11901_/CLK line[105] VGND VGND VPWR VPWR _11903_/Q sky130_fd_sc_hd__dfxtp_1
X_12883_ _12881_/CLK line[41] VGND VGND VPWR VPWR _12883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11834_ _11833_/Q _11837_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_11765_ _11765_/CLK _11766_/X VGND VGND VPWR VPWR _11757_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11840__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[22\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _13932_/X wr VGND VGND VPWR VPWR _10716_/X sky130_fd_sc_hd__and2_1
X_13504_ _13503_/Q _13517_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11872_/A wr VGND VGND VPWR VPWR _11696_/X sky130_fd_sc_hd__and2_1
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10456__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10647_ _13932_/X VGND VGND VPWR VPWR _10647_/Y sky130_fd_sc_hd__inv_2
X_13435_ _13439_/CLK line[37] VGND VGND VPWR VPWR _13436_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].CGAND_A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[19\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13365_/Q _13377_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_10578_ _10594_/CLK line[16] VGND VGND VPWR VPWR _10579_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13767__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12671__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12317_ _12311_/CLK line[38] VGND VGND VPWR VPWR _12317_/Q sky130_fd_sc_hd__dfxtp_1
X_13297_ _13285_/CLK line[102] VGND VGND VPWR VPWR _13297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07765__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12248_ _12247_/Q _12257_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_12179_ _12177_/CLK line[103] VGND VGND VPWR VPWR _12180_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[21\].VALID\[8\].FF OVHB\[21\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[21\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06740_ _06740_/CLK line[63] VGND VGND VPWR VPWR _06740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06671_ _06670_/Q _06692_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13007__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08410_ _08410_/CLK line[58] VGND VGND VPWR VPWR _08411_/A sky130_fd_sc_hd__dfxtp_1
X_05622_ _05632_/CLK line[49] VGND VGND VPWR VPWR _05623_/A sky130_fd_sc_hd__dfxtp_1
X_09390_ _09414_/CLK line[122] VGND VGND VPWR VPWR _09390_/Q sky130_fd_sc_hd__dfxtp_1
X_08341_ _08341_/A _08372_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12846__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05553_ _05553_/A _05572_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[21\].VALID\[5\].TOBUF OVHB\[21\].VALID\[5\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[29\].CG clk OVHB\[29\].CGAND/X VGND VGND VPWR VPWR OVHB\[29\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_71_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08272_ _08282_/CLK line[123] VGND VGND VPWR VPWR _08272_/Q sky130_fd_sc_hd__dfxtp_1
X_05484_ _05476_/CLK line[114] VGND VGND VPWR VPWR _05484_/Q sky130_fd_sc_hd__dfxtp_1
X_07223_ _07222_/Q _07252_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07154_ _07170_/CLK line[124] VGND VGND VPWR VPWR _07155_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06105_ _06104_/Q _06132_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12581__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07085_ _07085_/A _07112_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07675__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06036_ _06050_/CLK line[125] VGND VGND VPWR VPWR _06036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11197__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09890__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07987_ _13920_/X VGND VGND VPWR VPWR _07987_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09726_ _09725_/Q _09737_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_06938_ _06960_/CLK line[16] VGND VGND VPWR VPWR _06938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05923__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09657_ _09659_/CLK line[102] VGND VGND VPWR VPWR _09657_/Q sky130_fd_sc_hd__dfxtp_1
X_06869_ _06869_/A _06902_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08608_ _08607_/Q _08617_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
X_09588_ _09587_/Q _09597_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[11\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08541_/CLK line[103] VGND VGND VPWR VPWR _08539_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12756__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06754__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _11549_/Q _11557_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09130__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ _10473_/CLK line[104] VGND VGND VPWR VPWR _10501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ _11479_/CLK line[40] VGND VGND VPWR VPWR _11482_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13220_ _13219_/Q _13237_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
X_10432_ _10431_/Q _10437_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13151_ _13163_/CLK line[35] VGND VGND VPWR VPWR _13152_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10363_ _10341_/CLK line[41] VGND VGND VPWR VPWR _10363_/Q sky130_fd_sc_hd__dfxtp_1
X_12102_ _12102_/A _12117_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[11\].TOBUF OVHB\[17\].VALID\[11\].FF/Q OVHB\[17\].INV/Y VGND VGND
+ VPWR VPWR _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13082_ _13081_/Q _13097_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_10294_ _10294_/A _10297_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12033_ _12019_/CLK line[36] VGND VGND VPWR VPWR _12033_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[7\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06929__D line[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13984_ _13982_/X _13990_/B _13990_/A _13990_/D VGND VGND VPWR VPWR _13984_/X sky130_fd_sc_hd__and4bb_4
XFILLER_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09305__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12935_ _12937_/CLK line[79] VGND VGND VPWR VPWR _12935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12866_ _12865_/Q _12887_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11817_ _11823_/CLK line[65] VGND VGND VPWR VPWR _11817_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11570__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12797_ _12803_/CLK line[1] VGND VGND VPWR VPWR _12797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06664__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11748_ _11747_/Q _11767_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09040__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[10\].TOBUF OVHB\[10\].VALID\[10\].FF/Q OVHB\[10\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10186__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ _11691_/CLK line[2] VGND VGND VPWR VPWR _11679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[15\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13418_ _13417_/Q _13447_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13497__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13349_ _13347_/CLK line[12] VGND VGND VPWR VPWR _13349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_MUX.MUX\[24\]_A0 _10887_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07910_ _07909_/Q _07917_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
X_08890_ _08889_/Q _08897_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07841_ _07837_/CLK line[40] VGND VGND VPWR VPWR _07842_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11745__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06839__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07772_ _07772_/A _07777_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_04984_ _05000_/CLK line[28] VGND VGND VPWR VPWR _04984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05743__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06201__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09215__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06723_ _06711_/CLK line[41] VGND VGND VPWR VPWR _06723_/Q sky130_fd_sc_hd__dfxtp_1
X_09511_ _09507_/CLK line[35] VGND VGND VPWR VPWR _09511_/Q sky130_fd_sc_hd__dfxtp_1
X_09442_ _09441_/Q _09457_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
X_06654_ _06653_/Q _06657_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05605_ _05605_/CLK _05606_/X VGND VGND VPWR VPWR _05575_/CLK sky130_fd_sc_hd__dlclkp_1
X_09373_ _09365_/CLK line[100] VGND VGND VPWR VPWR _09373_/Q sky130_fd_sc_hd__dfxtp_1
X_06585_ _06585_/CLK _06586_/X VGND VGND VPWR VPWR _06565_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_127_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08324_ _08323_/Q _08337_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_05536_ _13909_/X wr VGND VGND VPWR VPWR _05536_/X sky130_fd_sc_hd__and2_1
XANTENNA__10096__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08255_ _08257_/CLK line[101] VGND VGND VPWR VPWR _08255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05467_ _13908_/X VGND VGND VPWR VPWR _05467_/Y sky130_fd_sc_hd__inv_2
X_07206_ _07205_/Q _07217_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[13\].FF_D A[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08186_ _08185_/Q _08197_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_05398_ _05424_/CLK line[80] VGND VGND VPWR VPWR _05398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07137_ _07117_/CLK line[102] VGND VGND VPWR VPWR _07137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05918__D line[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07068_ _07067_/Q _07077_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06019_ _06023_/CLK line[103] VGND VGND VPWR VPWR _06020_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05653__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[10\].TOBUF OVHB\[30\].VALID\[10\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
X_09709_ _09721_/CLK line[12] VGND VGND VPWR VPWR _09709_/Q sky130_fd_sc_hd__dfxtp_1
X_10981_ _10977_/CLK line[67] VGND VGND VPWR VPWR _10982_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13870__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[25\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12720_ _12720_/A _12747_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12486__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _12667_/CLK line[77] VGND VGND VPWR VPWR _12652_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11601_/Q _11627_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12581_/Q _12607_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[3\].VALID\[2\].TOBUF OVHB\[3\].VALID\[2\].FF/Q OVHB\[3\].INV/Y VGND VGND VPWR
+ VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[28\].VALID\[8\].FF_D A[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _11535_/CLK line[78] VGND VGND VPWR VPWR _11534_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[5\].TOBUF OVHB\[28\].VALID\[5\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04937_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09795__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _11463_/Q _11487_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_13203_ _13213_/CLK line[64] VGND VGND VPWR VPWR _13203_/Q sky130_fd_sc_hd__dfxtp_1
X_10415_ _10405_/CLK line[79] VGND VGND VPWR VPWR _10415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10734__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11395_ _11395_/CLK line[15] VGND VGND VPWR VPWR _11395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13110__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05828__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[27\].VOBUF OVHB\[27\].V/Q OVHB\[27\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_10346_ _10345_/Q _10367_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
X_13134_ _13133_/Q _13167_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[9\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _13690_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08204__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13065_ _13075_/CLK line[10] VGND VGND VPWR VPWR _13066_/A sky130_fd_sc_hd__dfxtp_1
X_10277_ _10277_/CLK line[1] VGND VGND VPWR VPWR _10277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12016_ _12015_/Q _12047_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _13958_/X _13964_/B _13960_/X _13966_/D VGND VGND VPWR VPWR _13967_/X sky130_fd_sc_hd__and4b_4
X_12918_ _12902_/CLK line[57] VGND VGND VPWR VPWR _12918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13898_ _13882_/CLK line[121] VGND VGND VPWR VPWR _13898_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10909__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12849_ _12848_/Q _12852_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06394__D line[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06370_ _06369_/Q _06377_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06972__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05321_ _05299_/CLK line[40] VGND VGND VPWR VPWR _05321_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[29\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _11030_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06691__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08040_ _08039_/Q _08057_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_05252_ _05252_/A _05257_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
X_05183_ _05157_/CLK line[105] VGND VGND VPWR VPWR _05183_/Q sky130_fd_sc_hd__dfxtp_1
X_09991_ _10011_/CLK line[13] VGND VGND VPWR VPWR _09992_/A sky130_fd_sc_hd__dfxtp_1
X_08942_ _08941_/Q _08967_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07953__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08873_ _08869_/CLK line[14] VGND VGND VPWR VPWR _08873_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11475__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07824_ _07823_/Q _07847_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06569__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07755_ _07773_/CLK line[15] VGND VGND VPWR VPWR _07756_/A sky130_fd_sc_hd__dfxtp_1
X_04967_ _04947_/CLK line[6] VGND VGND VPWR VPWR _04967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06866__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06706_ _06706_/A _06727_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08784__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07686_ _07686_/A _07707_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06637_ _06633_/CLK line[1] VGND VGND VPWR VPWR _06637_/Q sky130_fd_sc_hd__dfxtp_1
X_09425_ _09427_/CLK line[10] VGND VGND VPWR VPWR _09426_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ _09356_/A _09387_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_06568_ _06568_/A _06587_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08307_ _08329_/CLK line[11] VGND VGND VPWR VPWR _08307_/Q sky130_fd_sc_hd__dfxtp_1
X_05519_ _05519_/CLK line[2] VGND VGND VPWR VPWR _05519_/Q sky130_fd_sc_hd__dfxtp_1
X_09287_ _09307_/CLK line[75] VGND VGND VPWR VPWR _09288_/A sky130_fd_sc_hd__dfxtp_1
X_06499_ _06489_/CLK line[66] VGND VGND VPWR VPWR _06499_/Q sky130_fd_sc_hd__dfxtp_1
X_08238_ _08237_/Q _08267_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08169_ _08175_/CLK line[76] VGND VGND VPWR VPWR _08169_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[6\].FF OVHB\[9\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[9\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10200_ _10199_/Q _10227_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[28\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _10645_/CLK sky130_fd_sc_hd__clkbuf_4
X_11180_ _11180_/A _11207_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
X_10131_ _10145_/CLK line[77] VGND VGND VPWR VPWR _10131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08959__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10062_ _10061_/Q _10087_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11385__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[7\].TOBUF OVHB\[1\].VALID\[7\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_125_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05383__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13821_ _13821_/A _13832_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[6\]_A0 _09448_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08694__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13752_ _13746_/CLK line[54] VGND VGND VPWR VPWR _13752_/Q sky130_fd_sc_hd__dfxtp_1
X_10964_ _10963_/Q _10997_/Y VGND VGND VPWR VPWR _05084_/Z sky130_fd_sc_hd__ebufn_2
X_12703_ _12702_/Q _12712_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13683_ _13682_/Q _13692_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
X_10895_ _10903_/CLK line[42] VGND VGND VPWR VPWR _10895_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _12638_/CLK line[55] VGND VGND VPWR VPWR _12634_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[23\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12564_/Q _12572_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _11500_/CLK line[56] VGND VGND VPWR VPWR _11516_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06942__D line[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12490_/CLK line[120] VGND VGND VPWR VPWR _12496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10464__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11447_ _11447_/A _11452_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05558__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11378_ _11370_/CLK line[121] VGND VGND VPWR VPWR _11378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08512__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13775__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13117_ _13116_/Q _13132_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_10329_ _10328_/Q _10332_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08869__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07773__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08231__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13048_ _13050_/CLK line[116] VGND VGND VPWR VPWR _13048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[21\]_A3 _07171_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[8\].FF OVHB\[7\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[7\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05870_ _05869_/Q _05887_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05293__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDATA\[17\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _07390_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07540_ _07539_/Q _07567_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10639__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07471_ _07467_/CLK line[13] VGND VGND VPWR VPWR _07471_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13015__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06422_ _06422_/A _06447_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_09210_ _09210_/CLK _09211_/X VGND VGND VPWR VPWR _09200_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08109__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09141_ _13923_/X wr VGND VGND VPWR VPWR _09141_/X sky130_fd_sc_hd__and2_1
XOVHB\[7\].V OVHB\[7\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[7\].V/Q sky130_fd_sc_hd__dfrtp_1
X_06353_ _06353_/CLK line[14] VGND VGND VPWR VPWR _06354_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08406__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07948__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05304_ _05303_/Q _05327_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09072_ _13923_/X VGND VGND VPWR VPWR _09072_/Y sky130_fd_sc_hd__inv_2
X_06284_ _06283_/Q _06307_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
X_08023_ _08033_/CLK line[0] VGND VGND VPWR VPWR _08023_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10374__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05235_ _05253_/CLK line[15] VGND VGND VPWR VPWR _05236_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[13\].TOBUF OVHB\[7\].VALID\[13\].FF/Q OVHB\[7\].INV/Y VGND VGND
+ VPWR VPWR _04920_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_128_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05468__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05166_ _05166_/A _05187_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
X_09974_ _09978_/CLK line[119] VGND VGND VPWR VPWR _09974_/Q sky130_fd_sc_hd__dfxtp_1
X_05097_ _05093_/CLK line[65] VGND VGND VPWR VPWR _05097_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07683__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08925_ _08924_/Q _08932_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06299__D line[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08856_ _08850_/CLK line[120] VGND VGND VPWR VPWR _08857_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[30\].V OVHB\[30\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[30\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05781__A _13909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07807_ _07806_/Q _07812_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05999_ _06023_/CLK line[108] VGND VGND VPWR VPWR _06000_/A sky130_fd_sc_hd__dfxtp_1
X_08787_ _08787_/A _08792_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07738_ _07724_/CLK line[121] VGND VGND VPWR VPWR _07739_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04932__B2 _04932_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05931__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__10549__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _07005_/CLK sky130_fd_sc_hd__clkbuf_4
X_07669_ _07668_/Q _07672_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09408_ _09414_/CLK line[116] VGND VGND VPWR VPWR _09409_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[12\].TOBUF OVHB\[0\].VALID\[12\].FF/Q OVHB\[0\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_10680_ _10680_/CLK _10681_/X VGND VGND VPWR VPWR _10656_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12764__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09339_ _09338_/Q _09352_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07858__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _12352_/CLK line[53] VGND VGND VPWR VPWR _12350_/Q sky130_fd_sc_hd__dfxtp_1
X_11301_ _11301_/A _11312_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_12281_ _12281_/A _12292_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11232_ _11216_/CLK line[54] VGND VGND VPWR VPWR _11232_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05956__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XOVHB\[23\].VALID\[13\].FF OVHB\[23\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[23\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11163_ _11162_/Q _11172_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10114_ _10100_/CLK line[55] VGND VGND VPWR VPWR _10114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11094_ _11090_/CLK line[119] VGND VGND VPWR VPWR _11094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12004__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10045_ _10044_/Q _10052_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[21\].V OVHB\[21\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[21\].V/Q sky130_fd_sc_hd__dfrtp_1
XOVHB\[16\].VALID\[0\].FF OVHB\[16\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[16\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12939__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13804_ _13822_/CLK line[92] VGND VGND VPWR VPWR _13805_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09313__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11996_ _12002_/CLK line[19] VGND VGND VPWR VPWR _11996_/Q sky130_fd_sc_hd__dfxtp_1
X_13735_ _13734_/Q _13762_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
X_10947_ _10947_/A _10962_/Y VGND VGND VPWR VPWR _10387_/Z sky130_fd_sc_hd__ebufn_2
X_13666_ _13682_/CLK line[29] VGND VGND VPWR VPWR _13666_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10878_ _10872_/CLK line[20] VGND VGND VPWR VPWR _10878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ _12616_/Q _12642_/Y VGND VGND VPWR VPWR _10377_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ _13596_/Q _13622_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06672__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12548_ _12560_/CLK line[30] VGND VGND VPWR VPWR _12548_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06027__A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12479_ _12478_/Q _12502_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09983__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05288__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05020_ _05019_/Q _05047_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[21\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08599__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06971_ _07111_/A wr VGND VGND VPWR VPWR _06971_/X sky130_fd_sc_hd__and2_1
XFILLER_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08896__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08710_ _08710_/CLK line[53] VGND VGND VPWR VPWR _08711_/A sky130_fd_sc_hd__dfxtp_1
X_05922_ _13910_/X VGND VGND VPWR VPWR _05922_/Y sky130_fd_sc_hd__inv_2
X_09690_ _09694_/CLK line[117] VGND VGND VPWR VPWR _09691_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].V OVHB\[12\].V/CLK TIE/HI rst_n VGND VGND VPWR VPWR OVHB\[12\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07008__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05853_ _05871_/CLK line[32] VGND VGND VPWR VPWR _05853_/Q sky130_fd_sc_hd__dfxtp_1
X_08641_ _08640_/Q _08652_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[7\].TOBUF OVHB\[8\].VALID\[7\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11753__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06847__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05784_ _05783_/Q _05817_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_08572_ _08560_/CLK line[118] VGND VGND VPWR VPWR _08572_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09223__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07523_ _07523_/A _07532_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07454_ _07446_/CLK line[119] VGND VGND VPWR VPWR _07455_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[2\].FF OVHB\[14\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[14\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07321__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06405_ _06404_/Q _06412_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07385_ _07385_/A _07392_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[31\].VALID\[6\].FF OVHB\[31\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[31\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09124_ _09116_/CLK line[114] VGND VGND VPWR VPWR _09124_/Q sky130_fd_sc_hd__dfxtp_1
X_06336_ _06320_/CLK line[120] VGND VGND VPWR VPWR _06336_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[14\].TOBUF OVHB\[23\].VALID\[14\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09055_ _09054_/Q _09072_/Y VGND VGND VPWR VPWR _07095_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06267_ _06266_/Q _06272_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10682__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05198__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08006_ _08000_/CLK line[115] VGND VGND VPWR VPWR _08007_/A sky130_fd_sc_hd__dfxtp_1
X_05218_ _05214_/CLK line[121] VGND VGND VPWR VPWR _05218_/Q sky130_fd_sc_hd__dfxtp_1
X_06198_ _06186_/CLK line[57] VGND VGND VPWR VPWR _06198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11928__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05149_ _05148_/Q _05152_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09957_ _09956_/Q _09982_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08908_ _08922_/CLK line[30] VGND VGND VPWR VPWR _08908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09888_ _09908_/CLK line[94] VGND VGND VPWR VPWR _09888_/Q sky130_fd_sc_hd__dfxtp_1
X_08839_ _08838_/Q _08862_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11663__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11850_ _11846_/CLK line[95] VGND VGND VPWR VPWR _11850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05661__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10801_ _10801_/A _10822_/Y VGND VGND VPWR VPWR _13601_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10279__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[3\]_A3 _13572_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11781_ _11781_/A _11802_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10857__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13520_ _13528_/CLK line[90] VGND VGND VPWR VPWR _13520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08972__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10732_ _10728_/CLK line[81] VGND VGND VPWR VPWR _10732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10576__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13451_ _13450_/Q _13482_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12494__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10663_ _10662_/Q _10682_/Y VGND VGND VPWR VPWR _07023_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[11\]_A2 _13488_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[2\].TOBUF OVHB\[15\].VALID\[2\].FF/Q OVHB\[15\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07588__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12402_ _12414_/CLK line[91] VGND VGND VPWR VPWR _12402_/Q sky130_fd_sc_hd__dfxtp_1
X_10594_ _10594_/CLK line[18] VGND VGND VPWR VPWR _10595_/A sky130_fd_sc_hd__dfxtp_1
X_13382_ _13394_/CLK line[27] VGND VGND VPWR VPWR _13383_/A sky130_fd_sc_hd__dfxtp_1
X_12333_ _12332_/Q _12362_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[12\].VALID\[4\].FF OVHB\[12\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[12\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12264_ _12268_/CLK line[28] VGND VGND VPWR VPWR _12264_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11838__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11215_ _11214_/Q _11242_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10742__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12195_ _12194_/Q _12222_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05836__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08212__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11146_ _11148_/CLK line[29] VGND VGND VPWR VPWR _11146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11077_ _11076_/Q _11102_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10028_ _10042_/CLK line[30] VGND VGND VPWR VPWR _10029_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12669__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11979_ _11978_/Q _12012_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09978__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13718_ _13717_/Q _13727_/Y VGND VGND VPWR VPWR _05038_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10917__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13649_ _13631_/CLK line[7] VGND VGND VPWR VPWR _13650_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07498__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07170_ _07170_/CLK line[117] VGND VGND VPWR VPWR _07170_/Q sky130_fd_sc_hd__dfxtp_1
X_06121_ _06120_/Q _06132_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
X_06052_ _06050_/CLK line[118] VGND VGND VPWR VPWR _06052_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[9\].FF OVHB\[28\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[28\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05003_ _05002_/Q _05012_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10652__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[1\].TOBUF OVHB\[21\].VALID\[1\].FF/Q OVHB\[21\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_09811_ _09810_/Q _09842_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09742_ _09760_/CLK line[27] VGND VGND VPWR VPWR _09742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12222__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06954_ _06960_/CLK line[18] VGND VGND VPWR VPWR _06955_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[6\].FF OVHB\[10\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[10\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07961__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12579__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05905_ _05904_/Q _05922_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
X_09673_ _09672_/Q _09702_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11483__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06885_ _06884_/Q _06902_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06577__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08624_ _08646_/CLK line[28] VGND VGND VPWR VPWR _08624_/Q sky130_fd_sc_hd__dfxtp_1
X_05836_ _05836_/CLK line[19] VGND VGND VPWR VPWR _05836_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[11\].INV _13953_/X VGND VGND VPWR VPWR OVHB\[11\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08554_/Q _08582_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
X_05767_ _05767_/A _05782_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09888__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07506_ _07518_/CLK line[29] VGND VGND VPWR VPWR _07507_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08486_ _08480_/CLK line[93] VGND VGND VPWR VPWR _08487_/A sky130_fd_sc_hd__dfxtp_1
X_05698_ _05708_/CLK line[84] VGND VGND VPWR VPWR _05698_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07437_ _07436_/Q _07462_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10827__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[26\].INV _13974_/X VGND VGND VPWR VPWR OVHB\[26\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_11_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__D line[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07986__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07368_ _07380_/CLK line[94] VGND VGND VPWR VPWR _07369_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07201__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09107_ _13923_/X VGND VGND VPWR VPWR _09107_/Y sky130_fd_sc_hd__inv_2
X_06319_ _06319_/A _06342_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
X_07299_ _07298_/Q _07322_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09038_ _09068_/CLK line[80] VGND VGND VPWR VPWR _09038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12116__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11658__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09128__D line[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11000_ _11002_/CLK line[90] VGND VGND VPWR VPWR _11000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOVHB\[13\].VALID\[7\].TOBUF OVHB\[13\].VALID\[7\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_12951_ _12937_/CLK line[72] VGND VGND VPWR VPWR _12951_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11393__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _11902_/A _11907_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06487__D line[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12882_ _12881_/Q _12887_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05391__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDATA\[7\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _13305_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11833_ _11823_/CLK line[73] VGND VGND VPWR VPWR _11833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11764_ _11763_/Q _11767_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08057__A _13940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13497_/CLK line[68] VGND VGND VPWR VPWR _13503_/Q sky130_fd_sc_hd__dfxtp_1
X_10715_ _10715_/CLK _10716_/X VGND VGND VPWR VPWR _10707_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_92_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11695_/CLK _11696_/X VGND VGND VPWR VPWR _11691_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13433_/Q _13447_/Y VGND VGND VPWR VPWR _05594_/Z sky130_fd_sc_hd__ebufn_2
X_10646_ _13932_/X wr VGND VGND VPWR VPWR _10646_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[26\].CGAND_B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[19\]_S1 A[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13365_ _13347_/CLK line[5] VGND VGND VPWR VPWR _13365_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10577_ _13932_/X VGND VGND VPWR VPWR _10577_/Y sky130_fd_sc_hd__inv_2
X_12316_ _12316_/A _12327_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06950__D line[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13296_ _13295_/Q _13307_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11568__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12247_ _12227_/CLK line[6] VGND VGND VPWR VPWR _12247_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05566__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09038__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12178_ _12178_/A _12187_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13783__D line[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08877__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11129_ _11111_/CLK line[7] VGND VGND VPWR VPWR _11130_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06670_ _06682_/CLK line[31] VGND VGND VPWR VPWR _06670_/Q sky130_fd_sc_hd__dfxtp_1
X_05621_ _05620_/Q _05642_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09351__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08340_ _08358_/CLK line[26] VGND VGND VPWR VPWR _08341_/A sky130_fd_sc_hd__dfxtp_1
X_05552_ _05568_/CLK line[17] VGND VGND VPWR VPWR _05553_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09501__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[6\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _12920_/CLK sky130_fd_sc_hd__clkbuf_4
X_08271_ _08270_/Q _08302_/Y VGND VGND VPWR VPWR _13591_/Z sky130_fd_sc_hd__ebufn_2
X_05483_ _05483_/A _05502_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13023__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07222_ _07232_/CLK line[27] VGND VGND VPWR VPWR _07222_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08117__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07153_ _07152_/Q _07182_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
X_06104_ _06108_/CLK line[28] VGND VGND VPWR VPWR _06104_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[23\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07084_ _07098_/CLK line[92] VGND VGND VPWR VPWR _07085_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10382__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06035_ _06034_/Q _06062_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__05476__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09526__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13693__D line[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[16\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07691__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07986_ _13920_/X wr VGND VGND VPWR VPWR _07986_/X sky130_fd_sc_hd__and2_1
XFILLER_75_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09725_ _09721_/CLK line[5] VGND VGND VPWR VPWR _09725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06937_ _07111_/A VGND VGND VPWR VPWR _06937_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12887__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09656_ _09655_/Q _09667_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _10260_/CLK sky130_fd_sc_hd__clkbuf_4
X_06868_ _06892_/CLK line[112] VGND VGND VPWR VPWR _06869_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08607_ _08609_/CLK line[6] VGND VGND VPWR VPWR _08607_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06100__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05819_ _05818_/Q _05852_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09587_ _09577_/CLK line[70] VGND VGND VPWR VPWR _09587_/Q sky130_fd_sc_hd__dfxtp_1
X_06799_ _06798_/Q _06832_/Y VGND VGND VPWR VPWR _05119_/Z sky130_fd_sc_hd__ebufn_2
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08537_/Q _08547_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10557__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _08473_/CLK line[71] VGND VGND VPWR VPWR _08469_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.MUX\[28\] _10865_/Z _07015_/Z _06525_/Z _13595_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[28] sky130_fd_sc_hd__mux4_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[12\].TOBUF OVHB\[13\].VALID\[12\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
X_10500_ _10499_/Q _10507_/Y VGND VGND VPWR VPWR _07140_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08027__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[13\].FF OVHB\[28\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[28\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11480_ _11479_/Q _11487_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13868__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10431_ _10405_/CLK line[72] VGND VGND VPWR VPWR _10431_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12772__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[5\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _12535_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07866__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11031__A _11032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13150_ _13149_/Q _13167_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10362_ _10361_/Q _10367_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
X_12101_ _12109_/CLK line[67] VGND VGND VPWR VPWR _12102_/A sky130_fd_sc_hd__dfxtp_1
X_13081_ _13075_/CLK line[3] VGND VGND VPWR VPWR _13081_/Q sky130_fd_sc_hd__dfxtp_1
X_10293_ _10277_/CLK line[9] VGND VGND VPWR VPWR _10294_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12032_ _12031_/Q _12047_/Y VGND VGND VPWR VPWR _05592_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[28\].VALID\[1\].TOBUF OVHB\[28\].VALID\[1\].FF/Q OVHB\[28\].INV/Y VGND VGND
+ VPWR VPWR _04938_/B2 sky130_fd_sc_hd__ebufn_2
X_13983_ _13990_/A _13990_/B _13982_/X _13990_/D VGND VGND VPWR VPWR _13983_/Y sky130_fd_sc_hd__nor4b_4
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13108__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ _12933_/Q _12957_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07106__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12947__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[23\].VOBUF OVHB\[23\].V/Q OVHB\[23\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_12865_ _12881_/CLK line[47] VGND VGND VPWR VPWR _12865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11206__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11816_ _11815_/Q _11837_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12796_ _12795_/Q _12817_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[25\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _09875_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[1\].VALID\[1\].FF OVHB\[1\].V/CLK A[10] VGND VGND VPWR VPWR OVHB\[1\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11747_ _11757_/CLK line[33] VGND VGND VPWR VPWR _11747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _11677_/Q _11697_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
X_13417_ _13439_/CLK line[43] VGND VGND VPWR VPWR _13417_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12682__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10629_ _10627_/CLK line[34] VGND VGND VPWR VPWR _10629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06680__D line[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13348_ _13347_/Q _13377_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11298__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13279_ _13285_/CLK line[108] VGND VGND VPWR VPWR _13279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09991__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[24\]_A1 _13477_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[6\].FF_D A[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10930__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07840_ _07839_/Q _07847_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ _07773_/CLK line[8] VGND VGND VPWR VPWR _07772_/A sky130_fd_sc_hd__dfxtp_1
X_04983_ _04982_/Q _05012_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_09510_ _09509_/Q _09527_/Y VGND VGND VPWR VPWR _05030_/Z sky130_fd_sc_hd__ebufn_2
X_06722_ _06722_/A _06727_/Y VGND VGND VPWR VPWR _10922_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07016__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09441_ _09427_/CLK line[3] VGND VGND VPWR VPWR _09441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12857__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06653_ _06633_/CLK line[9] VGND VGND VPWR VPWR _06653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11761__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05604_ _05604_/A _05607_/Y VGND VGND VPWR VPWR _12884_/Z sky130_fd_sc_hd__ebufn_2
X_09372_ _09372_/A _09387_/Y VGND VGND VPWR VPWR _13572_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06855__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06584_ _06583_/Q _06587_/Y VGND VGND VPWR VPWR _06864_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09231__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08323_ _08329_/CLK line[4] VGND VGND VPWR VPWR _08323_/Q sky130_fd_sc_hd__dfxtp_1
X_05535_ _05535_/CLK _05536_/X VGND VGND VPWR VPWR _05519_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[12\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05466_ _13908_/X wr VGND VGND VPWR VPWR _05466_/X sky130_fd_sc_hd__and2_1
X_08254_ _08253_/Q _08267_/Y VGND VGND VPWR VPWR _06854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13688__D line[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07205_ _07183_/CLK line[5] VGND VGND VPWR VPWR _07205_/Q sky130_fd_sc_hd__dfxtp_1
X_05397_ _13908_/X VGND VGND VPWR VPWR _05397_/Y sky130_fd_sc_hd__inv_2
X_08185_ _08175_/CLK line[69] VGND VGND VPWR VPWR _08185_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _09490_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06590__D line[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07136_ _07135_/Q _07147_/Y VGND VGND VPWR VPWR _05176_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDATA\[14\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _06620_/CLK sky130_fd_sc_hd__clkbuf_4
X_07067_ _07043_/CLK line[70] VGND VGND VPWR VPWR _07067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06018_ _06017_/Q _06027_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11936__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09406__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[13\].FF OVHB\[0\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[0\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07969_ _07981_/CLK line[98] VGND VGND VPWR VPWR _07970_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09708_ _09708_/A _09737_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
X_10980_ _10979_/Q _10997_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[31\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09639_ _09659_/CLK line[108] VGND VGND VPWR VPWR _09639_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11671__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12649_/Q _12677_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06765__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _11605_/CLK line[109] VGND VGND VPWR VPWR _11601_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10287__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12601_/CLK line[45] VGND VGND VPWR VPWR _12581_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08980__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _11531_/Q _11557_/Y VGND VGND VPWR VPWR _10972_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[3\].TOBUF OVHB\[1\].VALID\[3\].FF/Q OVHB\[1\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13598__D line[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ _11479_/CLK line[46] VGND VGND VPWR VPWR _11463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[26\].VALID\[6\].TOBUF OVHB\[26\].VALID\[6\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__07596__D line[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13202_ _13272_/A VGND VGND VPWR VPWR _13202_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10414_ _10413_/Q _10437_/Y VGND VGND VPWR VPWR _13494_/Z sky130_fd_sc_hd__ebufn_2
X_11394_ _11393_/Q _11417_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
X_13133_ _13163_/CLK line[32] VGND VGND VPWR VPWR _13133_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11696__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10345_ _10341_/CLK line[47] VGND VGND VPWR VPWR _10345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06005__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13064_ _13063_/Q _13097_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_10276_ _10275_/Q _10297_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11846__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _12019_/CLK line[42] VGND VGND VPWR VPWR _12015_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].CG clk OVHB\[19\].CGAND/X VGND VGND VPWR VPWR OVHB\[19\].V/CLK sky130_fd_sc_hd__dlclkp_1
XDATA\[13\].CLKBUF\[4\] clk VGND VGND VPWR VPWR _06235_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_79_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__05844__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08220__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ _13964_/B _13958_/X _13960_/X _13966_/D VGND VGND VPWR VPWR _13966_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12917_ _12916_/Q _12922_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[24\].VALID\[11\].FF OVHB\[24\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[24\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13897_ _13897_/A _13902_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12848_ _12820_/CLK line[25] VGND VGND VPWR VPWR _12848_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10197__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12779_ _12778_/Q _12782_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
X_05320_ _05319_/Q _05327_/Y VGND VGND VPWR VPWR _05600_/Z sky130_fd_sc_hd__ebufn_2
X_05251_ _05253_/CLK line[8] VGND VGND VPWR VPWR _05252_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13301__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05182_ _05181_/Q _05187_/Y VGND VGND VPWR VPWR _13582_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09990_ _09989_/Q _10017_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[12\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08941_ _08947_/CLK line[45] VGND VGND VPWR VPWR _08941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[14\].VALID\[13\].FF OVHB\[14\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[14\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10660__D line[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08872_ _08871_/Q _08897_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05754__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07823_ _07837_/CLK line[46] VGND VGND VPWR VPWR _07823_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08130__D line[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07754_ _07753_/Q _07777_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04966_ _04965_/Q _04977_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[12\].CLKBUF\[1\] clk VGND VGND VPWR VPWR _05850_/CLK sky130_fd_sc_hd__clkbuf_4
X_06705_ _06711_/CLK line[47] VGND VGND VPWR VPWR _06706_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12587__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07685_ _07679_/CLK line[111] VGND VGND VPWR VPWR _07686_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09424_ _09423_/Q _09457_/Y VGND VGND VPWR VPWR _06904_/Z sky130_fd_sc_hd__ebufn_2
X_06636_ _06636_/A _06657_/Y VGND VGND VPWR VPWR _11396_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09355_ _09365_/CLK line[106] VGND VGND VPWR VPWR _09356_/A sky130_fd_sc_hd__dfxtp_1
X_06567_ _06565_/CLK line[97] VGND VGND VPWR VPWR _06568_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09896__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08306_ _08305_/Q _08337_/Y VGND VGND VPWR VPWR _11386_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13061__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05518_ _05517_/Q _05537_/Y VGND VGND VPWR VPWR _04958_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09286_ _09285_/Q _09317_/Y VGND VGND VPWR VPWR _13486_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06498_ _06497_/Q _06517_/Y VGND VGND VPWR VPWR _13498_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08237_ _08257_/CLK line[107] VGND VGND VPWR VPWR _08237_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10835__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05449_ _05445_/CLK line[98] VGND VGND VPWR VPWR _05449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13211__D line[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05929__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08305__D line[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08168_ _08167_/Q _08197_/Y VGND VGND VPWR VPWR _13488_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[10\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07119_ _07117_/CLK line[108] VGND VGND VPWR VPWR _07120_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08099_ _08113_/CLK line[44] VGND VGND VPWR VPWR _08100_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[24\].VALID\[0\].FF OVHB\[24\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[24\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10130_ _10129_/Q _10157_/Y VGND VGND VPWR VPWR _13490_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10061_ _10073_/CLK line[45] VGND VGND VPWR VPWR _10061_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09136__D line[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13236__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _13822_/CLK line[85] VGND VGND VPWR VPWR _13821_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[6\]_A1 _05038_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13751_ _13751_/A _13762_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
X_10963_ _10977_/CLK line[64] VGND VGND VPWR VPWR _10963_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].CGAND _11872_/A wr VGND VGND VPWR VPWR OVHB\[31\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA_DATA\[3\].CLKBUF\[3\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12702_ _12708_/CLK line[86] VGND VGND VPWR VPWR _12702_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06495__D line[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13682_ _13682_/CLK line[22] VGND VGND VPWR VPWR _13682_/Q sky130_fd_sc_hd__dfxtp_1
X_10894_ _10893_/Q _10927_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _12632_/Q _12642_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.MUX\[14\]_A0 _11394_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _12560_/CLK line[23] VGND VGND VPWR VPWR _12564_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11515_ _11514_/Q _11522_/Y VGND VGND VPWR VPWR _09555_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12494_/Q _12502_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11446_ _11440_/CLK line[24] VGND VGND VPWR VPWR _11447_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[25\].VALID\[9\].FF_D A[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12960__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11377_ _11377_/A _11382_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_13116_ _13120_/CLK line[19] VGND VGND VPWR VPWR _13116_/Q sky130_fd_sc_hd__dfxtp_1
X_10328_ _10314_/CLK line[25] VGND VGND VPWR VPWR _10328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11576__D line[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13047_ _13046_/Q _13062_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_10259_ _10259_/A _10262_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09046__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13791__D line[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08885__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[2\].FF OVHB\[22\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[22\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13949_ A_h[6] VGND VGND VPWR VPWR _13950_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__12200__D line[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07470_ _07469_/Q _07497_/Y VGND VGND VPWR VPWR _10830_/Z sky130_fd_sc_hd__ebufn_2
X_06421_ _06421_/CLK line[45] VGND VGND VPWR VPWR _06422_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[14\].TOBUF OVHB\[3\].VALID\[14\].FF/Q OVHB\[3\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XFILLER_72_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09140_ _09140_/CLK _09141_/X VGND VGND VPWR VPWR _09116_/CLK sky130_fd_sc_hd__dlclkp_1
X_06352_ _06351_/Q _06377_/Y VGND VGND VPWR VPWR _13352_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05303_ _05299_/CLK line[46] VGND VGND VPWR VPWR _05303_/Q sky130_fd_sc_hd__dfxtp_1
X_06283_ _06285_/CLK line[110] VGND VGND VPWR VPWR _06283_/Q sky130_fd_sc_hd__dfxtp_1
X_09071_ _13923_/X wr VGND VGND VPWR VPWR _09071_/X sky130_fd_sc_hd__and2_1
X_08022_ _13920_/X VGND VGND VPWR VPWR _08022_/Y sky130_fd_sc_hd__inv_2
XOVHB\[8\].VALID\[3\].TOBUF OVHB\[8\].VALID\[3\].FF/Q OVHB\[8\].INV/Y VGND VGND VPWR
+ VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
X_05234_ _05233_/Q _05257_/Y VGND VGND VPWR VPWR _11394_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[14\].FF_D A[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05165_ _05157_/CLK line[111] VGND VGND VPWR VPWR _05166_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09973_ _09973_/A _09982_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_05096_ _05095_/Q _05117_/Y VGND VGND VPWR VPWR _13496_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10390__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08924_ _08922_/CLK line[23] VGND VGND VPWR VPWR _08924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05484__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08855_ _08854_/Q _08862_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XOVHB\[23\].VALID\[10\].TOBUF OVHB\[23\].VALID\[10\].FF/Q OVHB\[23\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05781__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07806_ _07788_/CLK line[24] VGND VGND VPWR VPWR _07806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08795__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08786_ _08762_/CLK line[88] VGND VGND VPWR VPWR _08787_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05998_ _05997_/Q _06027_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
X_07737_ _07737_/A _07742_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_04949_ _04947_/CLK line[12] VGND VGND VPWR VPWR _04949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07668_ _07644_/CLK line[89] VGND VGND VPWR VPWR _07668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09407_ _09406_/Q _09422_/Y VGND VGND VPWR VPWR _07167_/Z sky130_fd_sc_hd__ebufn_2
X_06619_ _06619_/A _06622_/Y VGND VGND VPWR VPWR _07179_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07599_ _07598_/Q _07602_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XOVHB\[20\].VALID\[4\].FF OVHB\[20\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[20\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09338_ _09320_/CLK line[84] VGND VGND VPWR VPWR _09338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XMUX.MUX\[10\] _11386_/Z _05576_/Z _13486_/Z _07116_/Z A[2] A[3] VGND VGND VPWR VPWR
+ Do[10] sky130_fd_sc_hd__mux4_1
XANTENNA__10565__D line[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09269_ _09268_/Q _09282_/Y VGND VGND VPWR VPWR _13469_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05659__D line[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11300_ _11302_/CLK line[85] VGND VGND VPWR VPWR _11301_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[11\].FF OVHB\[10\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[10\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08035__D line[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12280_ _12268_/CLK line[21] VGND VGND VPWR VPWR _12281_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13876__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11231_ _11230_/Q _11242_/Y VGND VGND VPWR VPWR _10391_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05956__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07874__D line[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11162_ _11148_/CLK line[22] VGND VGND VPWR VPWR _11162_/Q sky130_fd_sc_hd__dfxtp_1
X_10113_ _10112_/Q _10122_/Y VGND VGND VPWR VPWR _13473_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11093_ _11092_/Q _11102_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
X_10044_ _10042_/CLK line[23] VGND VGND VPWR VPWR _10044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13803_ _13802_/Q _13832_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
X_11995_ _11994_/Q _12012_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13116__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13734_ _13746_/CLK line[60] VGND VGND VPWR VPWR _13734_/Q sky130_fd_sc_hd__dfxtp_1
X_10946_ _10930_/CLK line[51] VGND VGND VPWR VPWR _10947_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[10\].FF_D A[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[5\].FF OVHB\[19\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[19\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13665_ _13665_/A _13692_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
X_10877_ _10876_/Q _10892_/Y VGND VGND VPWR VPWR _10877_/Z sky130_fd_sc_hd__ebufn_2
X_12616_ _12638_/CLK line[61] VGND VGND VPWR VPWR _12616_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ _13598_/CLK line[125] VGND VGND VPWR VPWR _13596_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10475__D line[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12547_ _12546_/Q _12572_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[1\].CLKBUF\[5\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12478_ _12490_/CLK line[126] VGND VGND VPWR VPWR _12478_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12690__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11429_ _11428_/Q _11452_/Y VGND VGND VPWR VPWR _09469_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07784__D line[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06970_ _06970_/CLK _06971_/X VGND VGND VPWR VPWR _06960_/CLK sky130_fd_sc_hd__dlclkp_1
X_05921_ _13910_/X wr VGND VGND VPWR VPWR _05921_/X sky130_fd_sc_hd__and2_1
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08640_ _08646_/CLK line[21] VGND VGND VPWR VPWR _08640_/Q sky130_fd_sc_hd__dfxtp_1
X_05852_ _13910_/X VGND VGND VPWR VPWR _05852_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08571_ _08570_/Q _08582_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[6\].VALID\[8\].TOBUF OVHB\[6\].VALID\[8\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_05783_ _05799_/CLK line[0] VGND VGND VPWR VPWR _05783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ _07518_/CLK line[22] VGND VGND VPWR VPWR _07523_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07024__D line[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07602__A _07672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12865__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07453_ _07452_/Q _07462_/Y VGND VGND VPWR VPWR _13613_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07959__D line[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06404_ _06408_/CLK line[23] VGND VGND VPWR VPWR _06404_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07321__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06863__D line[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07384_ _07380_/CLK line[87] VGND VGND VPWR VPWR _07385_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09123_ _09122_/Q _09142_/Y VGND VGND VPWR VPWR _05203_/Z sky130_fd_sc_hd__ebufn_2
X_06335_ _06334_/Q _06342_/Y VGND VGND VPWR VPWR _09415_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09054_ _09068_/CLK line[82] VGND VGND VPWR VPWR _09054_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[7\].FF OVHB\[17\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[17\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06266_ _06244_/CLK line[88] VGND VGND VPWR VPWR _06266_/Q sky130_fd_sc_hd__dfxtp_1
X_08005_ _08004_/Q _08022_/Y VGND VGND VPWR VPWR _13605_/Z sky130_fd_sc_hd__ebufn_2
X_05217_ _05217_/A _05222_/Y VGND VGND VPWR VPWR _12777_/Z sky130_fd_sc_hd__ebufn_2
X_06197_ _06196_/Q _06202_/Y VGND VGND VPWR VPWR _13477_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[5\].VALID\[13\].FF OVHB\[5\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[5\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05148_ _05122_/CLK line[89] VGND VGND VPWR VPWR _05148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12105__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05079_ _05079_/A _05082_/Y VGND VGND VPWR VPWR _07039_/Z sky130_fd_sc_hd__ebufn_2
X_09956_ _09978_/CLK line[125] VGND VGND VPWR VPWR _09956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08907_ _08907_/A _08932_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09887_ _09887_/A _09912_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDATA\[3\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _12150_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08838_ _08850_/CLK line[126] VGND VGND VPWR VPWR _08838_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09414__D line[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08769_ _08768_/Q _08792_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
X_10800_ _10804_/CLK line[127] VGND VGND VPWR VPWR _10801_/A sky130_fd_sc_hd__dfxtp_1
X_11780_ _11776_/CLK line[63] VGND VGND VPWR VPWR _11781_/A sky130_fd_sc_hd__dfxtp_1
X_10731_ _10730_/Q _10752_/Y VGND VGND VPWR VPWR _11851_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13450_ _13468_/CLK line[58] VGND VGND VPWR VPWR _13450_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06773__D line[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10662_ _10656_/CLK line[49] VGND VGND VPWR VPWR _10662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_MUX.MUX\[11\]_A3 _07118_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12401_ _12400_/Q _12432_/Y VGND VGND VPWR VPWR _06521_/Z sky130_fd_sc_hd__ebufn_2
X_13381_ _13381_/A _13412_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_10593_ _10592_/Q _10612_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[3\].TOBUF OVHB\[13\].VALID\[3\].FF/Q OVHB\[13\].INV/Y VGND VGND
+ VPWR VPWR _04927_/A sky130_fd_sc_hd__ebufn_2
XANTENNA__05389__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12332_ _12352_/CLK line[59] VGND VGND VPWR VPWR _12332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12263_ _12263_/A _12292_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_11214_ _11216_/CLK line[60] VGND VGND VPWR VPWR _11214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12194_ _12204_/CLK line[124] VGND VGND VPWR VPWR _12194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12015__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11145_ _11144_/Q _11172_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[9\].FF OVHB\[15\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[15\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[11\].FF OVHB\[29\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[29\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06013__D line[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11076_ _11090_/CLK line[125] VGND VGND VPWR VPWR _11076_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11854__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10027_ _10026_/Q _10052_/Y VGND VGND VPWR VPWR _10867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06948__D line[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09324__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11978_ _12002_/CLK line[16] VGND VGND VPWR VPWR _11978_/Q sky130_fd_sc_hd__dfxtp_1
XDATA\[2\].CLKBUF\[2\] clk VGND VGND VPWR VPWR _11205_/CLK sky130_fd_sc_hd__clkbuf_4
X_13717_ _13701_/CLK line[38] VGND VGND VPWR VPWR _13717_/Q sky130_fd_sc_hd__dfxtp_1
X_10929_ _10928_/Q _10962_/Y VGND VGND VPWR VPWR _07009_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ _13648_/A _13657_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13579_ _13559_/CLK line[103] VGND VGND VPWR VPWR _13580_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].CG clk OVHB\[1\].CGAND/X VGND VGND VPWR VPWR OVHB\[1\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05299__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06120_ _06108_/CLK line[21] VGND VGND VPWR VPWR _06120_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[13\].FF OVHB\[19\].V/CLK A[22] VGND VGND VPWR VPWR OVHB\[19\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06051_ _06050_/Q _06062_/Y VGND VGND VPWR VPWR _07171_/Z sky130_fd_sc_hd__ebufn_2
X_05002_ _05000_/CLK line[22] VGND VGND VPWR VPWR _05002_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08403__D line[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[18\].VOBUF OVHB\[18\].V/Q OVHB\[18\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_09810_ _09834_/CLK line[58] VGND VGND VPWR VPWR _09810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09741_ _09740_/Q _09772_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_06953_ _06952_/Q _06972_/Y VGND VGND VPWR VPWR _10873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDATA\[22\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _09105_/CLK sky130_fd_sc_hd__clkbuf_4
X_05904_ _05902_/CLK line[50] VGND VGND VPWR VPWR _05904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09672_ _09694_/CLK line[123] VGND VGND VPWR VPWR _09672_/Q sky130_fd_sc_hd__dfxtp_1
X_06884_ _06892_/CLK line[114] VGND VGND VPWR VPWR _06884_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05762__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__05117__A _05152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08623_ _08622_/Q _08652_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05835_ _05835_/A _05852_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08560_/CLK line[124] VGND VGND VPWR VPWR _08554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05766_ _05756_/CLK line[115] VGND VGND VPWR VPWR _05767_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07505_ _07504_/Q _07532_/Y VGND VGND VPWR VPWR _10865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__D line[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08485_ _08485_/A _08512_/Y VGND VGND VPWR VPWR _06525_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05697_ _05697_/A _05712_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07689__D line[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07436_ _07446_/CLK line[125] VGND VGND VPWR VPWR _07436_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07986__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07367_ _07367_/A _07392_/Y VGND VGND VPWR VPWR _07087_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11004__D line[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09106_ _13923_/X wr VGND VGND VPWR VPWR _09106_/X sky130_fd_sc_hd__and2_1
X_06318_ _06320_/CLK line[126] VGND VGND VPWR VPWR _06319_/A sky130_fd_sc_hd__dfxtp_1
X_07298_ _07292_/CLK line[62] VGND VGND VPWR VPWR _07298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05002__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09037_ _13923_/X VGND VGND VPWR VPWR _09037_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10843__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06249_ _06248_/Q _06272_/Y VGND VGND VPWR VPWR _09609_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05937__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08313__D line[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09939_ _09925_/CLK line[103] VGND VGND VPWR VPWR _09939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06411__A _06551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[0\].FF_D A[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12950_ _12949_/Q _12957_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[11\].VALID\[8\].TOBUF OVHB\[11\].VALID\[8\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11901_ _11901_/CLK line[104] VGND VGND VPWR VPWR _11902_/A sky130_fd_sc_hd__dfxtp_1
X_12881_ _12881_/CLK line[40] VGND VGND VPWR VPWR _12881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11832_ _11831_/Q _11837_/Y VGND VGND VPWR VPWR _10992_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[21\].CLKBUF\[3\] clk VGND VGND VPWR VPWR _08720_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_42_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11763_ _11757_/CLK line[41] VGND VGND VPWR VPWR _11763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].VALID\[4\].FF_D A[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10713_/Q _10717_/Y VGND VGND VPWR VPWR _13514_/Z sky130_fd_sc_hd__ebufn_2
X_13502_ _13501_/Q _13517_/Y VGND VGND VPWR VPWR _13502_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11693_/Q _11697_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[11\].FF OVHB\[1\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[1\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13433_ _13439_/CLK line[36] VGND VGND VPWR VPWR _13433_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10645_ _10645_/CLK _10646_/X VGND VGND VPWR VPWR _10627_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_10_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13364_ _13363_/Q _13377_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10576_ _13932_/X wr VGND VGND VPWR VPWR _10576_/X sky130_fd_sc_hd__and2_1
XFILLER_10_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10753__D line[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12315_ _12311_/CLK line[37] VGND VGND VPWR VPWR _12316_/A sky130_fd_sc_hd__dfxtp_1
X_13295_ _13285_/CLK line[101] VGND VGND VPWR VPWR _13295_/Q sky130_fd_sc_hd__dfxtp_1
X_12246_ _12246_/A _12257_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12177_ _12177_/CLK line[102] VGND VGND VPWR VPWR _12178_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11128_ _11127_/Q _11137_/Y VGND VGND VPWR VPWR _09448_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11584__D line[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[2\].FF OVHB\[8\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[8\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].CG_CLK clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11059_ _11063_/CLK line[103] VGND VGND VPWR VPWR _11060_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06678__D line[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09054__D line[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09632__A _09632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[20\].CLKBUF\[1\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09989__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05620_ _05632_/CLK line[63] VGND VGND VPWR VPWR _05620_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08893__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09351__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10928__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05551_ _05550_/Q _05572_/Y VGND VGND VPWR VPWR _10871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08270_ _08282_/CLK line[122] VGND VGND VPWR VPWR _08270_/Q sky130_fd_sc_hd__dfxtp_1
X_05482_ _05476_/CLK line[113] VGND VGND VPWR VPWR _05483_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07302__D line[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[14\].TOBUF OVHB\[16\].VALID\[14\].FF/Q OVHB\[16\].INV/Y VGND VGND
+ VPWR VPWR _04923_/B sky130_fd_sc_hd__ebufn_2
XDATA\[20\].CLKBUF\[0\] clk VGND VGND VPWR VPWR _08335_/CLK sky130_fd_sc_hd__clkbuf_4
X_07221_ _07221_/A _07252_/Y VGND VGND VPWR VPWR _11421_/Z sky130_fd_sc_hd__ebufn_2
X_07152_ _07170_/CLK line[123] VGND VGND VPWR VPWR _07152_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[15\].VALID\[12\].FF_D A[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[6\] clk VGND VGND VPWR VPWR _05465_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_9_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11759__D line[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06103_ _06103_/A _06132_/Y VGND VGND VPWR VPWR _10863_/Z sky130_fd_sc_hd__ebufn_2
X_07083_ _07082_/Q _07112_/Y VGND VGND VPWR VPWR _11003_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09229__D line[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[1\]_S0 A[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06034_ _06050_/CLK line[124] VGND VGND VPWR VPWR _06034_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09807__A _09912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09526__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07985_ _07985_/CLK _07986_/X VGND VGND VPWR VPWR _07981_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11494__D line[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09724_ _09723_/Q _09737_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_06936_ _07111_/A wr VGND VGND VPWR VPWR _06936_/X sky130_fd_sc_hd__and2_1
XANTENNA__06588__D line[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__05492__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09655_ _09659_/CLK line[101] VGND VGND VPWR VPWR _09655_/Q sky130_fd_sc_hd__dfxtp_1
X_06867_ _06832_/A VGND VGND VPWR VPWR _06867_/Y sky130_fd_sc_hd__inv_2
X_08606_ _08606_/A _08617_/Y VGND VGND VPWR VPWR _10846_/Z sky130_fd_sc_hd__ebufn_2
X_05818_ _05836_/CLK line[16] VGND VGND VPWR VPWR _05818_/Q sky130_fd_sc_hd__dfxtp_1
X_09586_ _09585_/Q _09597_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
X_06798_ _06802_/CLK line[80] VGND VGND VPWR VPWR _06798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08541_/CLK line[102] VGND VGND VPWR VPWR _08537_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[4\].FF OVHB\[6\].V/CLK A[13] VGND VGND VPWR VPWR OVHB\[6\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05749_ _05748_/Q _05782_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[15\].VALID\[11\].FF OVHB\[15\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[15\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _08468_/A _08477_/Y VGND VGND VPWR VPWR _13508_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _07393_/CLK line[103] VGND VGND VPWR VPWR _07419_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ _08383_/CLK line[39] VGND VGND VPWR VPWR _08399_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].V_D TIE/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11312__A _11311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10430_ _10429_/Q _10437_/Y VGND VGND VPWR VPWR _13510_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11669__D line[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11031__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10573__D line[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10361_ _10341_/CLK line[40] VGND VGND VPWR VPWR _10361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__05667__D line[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12100_ _12100_/A _12117_/Y VGND VGND VPWR VPWR _06780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08043__D line[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13080_ _13079_/Q _13097_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_10292_ _10292_/A _10297_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13884__D line[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12031_ _12019_/CLK line[35] VGND VGND VPWR VPWR _12031_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08978__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[19\].CLKBUF\[2\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13982_ A_h[6] VGND VGND VPWR VPWR _13982_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[26\].VALID\[2\].TOBUF OVHB\[26\].VALID\[2\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12933_ _12937_/CLK line[78] VGND VGND VPWR VPWR _12933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12864_ _12864_/A _12887_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09602__D line[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11206__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11815_ _11823_/CLK line[79] VGND VGND VPWR VPWR _11815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10748__D line[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12795_ _12803_/CLK line[15] VGND VGND VPWR VPWR _12795_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13124__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11746_ _11746_/A _11767_/Y VGND VGND VPWR VPWR _05586_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08218__D line[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11691_/CLK line[1] VGND VGND VPWR VPWR _11677_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10628_ _10628_/A _10647_/Y VGND VGND VPWR VPWR _13428_/Z sky130_fd_sc_hd__ebufn_2
X_13416_ _13415_/Q _13447_/Y VGND VGND VPWR VPWR _05576_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[4\].VALID\[6\].FF OVHB\[4\].V/CLK A[15] VGND VGND VPWR VPWR OVHB\[4\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10483__D line[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13347_ _13347_/CLK line[11] VGND VGND VPWR VPWR _13347_/Q sky130_fd_sc_hd__dfxtp_1
X_10559_ _10571_/CLK line[2] VGND VGND VPWR VPWR _10559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05577__D line[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[10\].INV _13952_/X VGND VGND VPWR VPWR OVHB\[10\].INV/Y sky130_fd_sc_hd__inv_2
X_13278_ _13277_/Q _13307_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].CGAND _10192_/A wr VGND VGND VPWR VPWR OVHB\[26\].CGAND/X sky130_fd_sc_hd__and2_4
X_12229_ _12227_/CLK line[12] VGND VGND VPWR VPWR _12229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[24\]_A2 _13547_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07792__D line[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07147__A _07111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[25\].INV _13973_/X VGND VGND VPWR VPWR OVHB\[25\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07770_ _07770_/A _07777_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
X_04982_ _05000_/CLK line[27] VGND VGND VPWR VPWR _04982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06721_ _06711_/CLK line[40] VGND VGND VPWR VPWR _06722_/A sky130_fd_sc_hd__dfxtp_1
X_09440_ _09440_/A _09457_/Y VGND VGND VPWR VPWR _09160_/Z sky130_fd_sc_hd__ebufn_2
X_06652_ _06651_/Q _06657_/Y VGND VGND VPWR VPWR _09452_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[8\].TOBUF OVHB\[18\].VALID\[8\].FF/Q OVHB\[18\].INV/Y VGND VGND
+ VPWR VPWR _04935_/B2 sky130_fd_sc_hd__ebufn_2
X_05603_ _05575_/CLK line[41] VGND VGND VPWR VPWR _05604_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10658__D line[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09371_ _09365_/CLK line[99] VGND VGND VPWR VPWR _09372_/A sky130_fd_sc_hd__dfxtp_1
X_06583_ _06565_/CLK line[105] VGND VGND VPWR VPWR _06583_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13034__D line[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08322_ _08321_/Q _08337_/Y VGND VGND VPWR VPWR _11402_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08128__D line[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05534_ _05533_/Q _05537_/Y VGND VGND VPWR VPWR _11414_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07032__D line[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08253_ _08257_/CLK line[100] VGND VGND VPWR VPWR _08253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12873__D line[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05465_ _05465_/CLK _05466_/X VGND VGND VPWR VPWR _05445_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07967__D line[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07204_ _07203_/Q _07217_/Y VGND VGND VPWR VPWR _10844_/Z sky130_fd_sc_hd__ebufn_2
X_08184_ _08184_/A _08197_/Y VGND VGND VPWR VPWR _13504_/Z sky130_fd_sc_hd__ebufn_2
X_05396_ _13908_/X wr VGND VGND VPWR VPWR _05396_/X sky130_fd_sc_hd__and2_1
X_07135_ _07117_/CLK line[101] VGND VGND VPWR VPWR _07135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07066_ _07066_/A _07077_/Y VGND VGND VPWR VPWR _13506_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08441__A _13921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06017_ _06023_/CLK line[102] VGND VGND VPWR VPWR _06017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[12\].CGAND_A _13910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[20\].VALID\[3\].FF_D A[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[8\].FF OVHB\[2\].V/CLK A[17] VGND VGND VPWR VPWR OVHB\[2\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__D line[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12113__D line[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07968_ _07967_/Q _07987_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07207__D line[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09707_ _09721_/CLK line[11] VGND VGND VPWR VPWR _09708_/A sky130_fd_sc_hd__dfxtp_1
X_06919_ _06923_/CLK line[2] VGND VGND VPWR VPWR _06920_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07899_ _07905_/CLK line[66] VGND VGND VPWR VPWR _07900_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[13\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09638_ _09638_/A _09667_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09569_ _09577_/CLK line[76] VGND VGND VPWR VPWR _09570_/A sky130_fd_sc_hd__dfxtp_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _11600_/A _11627_/Y VGND VGND VPWR VPWR _06840_/Z sky130_fd_sc_hd__ebufn_2
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12580_/A _12607_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__A _13922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12783__D line[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11531_ _11535_/CLK line[77] VGND VGND VPWR VPWR _11531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06781__D line[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11462_ _11462_/A _11487_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11399__D line[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13201_ _13272_/A wr VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__and2_1
XANTENNA__11977__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10413_ _10405_/CLK line[78] VGND VGND VPWR VPWR _10413_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[7\].TOBUF OVHB\[24\].VALID\[7\].FF/Q OVHB\[24\].INV/Y VGND VGND
+ VPWR VPWR _04918_/A2 sky130_fd_sc_hd__ebufn_2
X_11393_ _11395_/CLK line[14] VGND VGND VPWR VPWR _11393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13132_ _13272_/A VGND VGND VPWR VPWR _13132_/Y sky130_fd_sc_hd__inv_2
X_10344_ _10343_/Q _10367_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11696__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13063_ _13075_/CLK line[0] VGND VGND VPWR VPWR _13063_/Q sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[2\].FF OVHB\[30\].V/CLK A[11] VGND VGND VPWR VPWR OVHB\[30\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10275_ _10277_/CLK line[15] VGND VGND VPWR VPWR _10275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12014_ _12013_/Q _12047_/Y VGND VGND VPWR VPWR _10894_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12023__D line[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07117__D line[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06021__D line[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12958__D line[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13965_ _13958_/X _13964_/B _13960_/X _13966_/D VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__11862__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12916_ _12902_/CLK line[56] VGND VGND VPWR VPWR _12916_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06956__D line[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10121__A _10192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13896_ _13882_/CLK line[120] VGND VGND VPWR VPWR _13897_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09332__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12847_ _12846_/Q _12852_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[17\].CLKBUF\[4\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12778_ _12774_/CLK line[121] VGND VGND VPWR VPWR _12778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13789__D line[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11729_ _11728_/Q _11732_/Y VGND VGND VPWR VPWR _10329_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05250_ _05249_/Q _05257_/Y VGND VGND VPWR VPWR _11410_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05181_ _05157_/CLK line[104] VGND VGND VPWR VPWR _05181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[29\].VALID\[3\].FF OVHB\[29\].V/CLK A[12] VGND VGND VPWR VPWR OVHB\[29\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08940_ _08940_/A _08967_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[10\].TOBUF OVHB\[3\].VALID\[10\].FF/Q OVHB\[3\].INV/Y VGND VGND
+ VPWR VPWR _04934_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09507__D line[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08871_ _08869_/CLK line[13] VGND VGND VPWR VPWR _08871_/Q sky130_fd_sc_hd__dfxtp_1
X_07822_ _07822_/A _07847_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[6\].TOBUF OVHB\[30\].VALID\[6\].FF/Q OVHB\[30\].INV/Y VGND VGND
+ VPWR VPWR _04924_/A sky130_fd_sc_hd__ebufn_2
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[0\].FF OVHB\[11\].V/CLK A[9] VGND VGND VPWR VPWR OVHB\[11\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[7\].FF_D A[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07753_ _07773_/CLK line[14] VGND VGND VPWR VPWR _07753_/Q sky130_fd_sc_hd__dfxtp_1
X_04965_ _04947_/CLK line[5] VGND VGND VPWR VPWR _04965_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11772__D line[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06704_ _06704_/A _06727_/Y VGND VGND VPWR VPWR _05584_/Z sky130_fd_sc_hd__ebufn_2
X_07684_ _07684_/A _07707_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05770__D line[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09423_ _09427_/CLK line[0] VGND VGND VPWR VPWR _09423_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10388__D line[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06635_ _06633_/CLK line[15] VGND VGND VPWR VPWR _06636_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13342__A _13272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09354_ _09353_/Q _09387_/Y VGND VGND VPWR VPWR _13554_/Z sky130_fd_sc_hd__ebufn_2
X_06566_ _06566_/A _06587_/Y VGND VGND VPWR VPWR _13566_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13699__D line[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08305_ _08329_/CLK line[10] VGND VGND VPWR VPWR _08305_/Q sky130_fd_sc_hd__dfxtp_1
X_05517_ _05519_/CLK line[1] VGND VGND VPWR VPWR _05517_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13061__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09285_ _09307_/CLK line[74] VGND VGND VPWR VPWR _09285_/Q sky130_fd_sc_hd__dfxtp_1
X_06497_ _06489_/CLK line[65] VGND VGND VPWR VPWR _06497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07697__D line[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08236_ _08235_/Q _08267_/Y VGND VGND VPWR VPWR _07116_/Z sky130_fd_sc_hd__ebufn_2
X_05448_ _05448_/A _05467_/Y VGND VGND VPWR VPWR _13568_/Z sky130_fd_sc_hd__ebufn_2
X_08167_ _08175_/CLK line[75] VGND VGND VPWR VPWR _08167_/Q sky130_fd_sc_hd__dfxtp_1
X_05379_ _05391_/CLK line[66] VGND VGND VPWR VPWR _05379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11012__D line[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07118_ _07117_/Q _07147_/Y VGND VGND VPWR VPWR _07118_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__06106__D line[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08098_ _08098_/A _08127_/Y VGND VGND VPWR VPWR _05578_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11947__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10851__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07049_ _07043_/CLK line[76] VGND VGND VPWR VPWR _07049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05945__D line[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10060_ _10059_/Q _10087_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08321__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13517__A _13552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XOVHB\[27\].VALID\[5\].FF OVHB\[27\].V/CLK A[14] VGND VGND VPWR VPWR OVHB\[27\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__04935__B1 A_h[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13236__B wr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12778__D line[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[6\]_A2 _13508_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[11\].FF OVHB\[6\].V/CLK A[20] VGND VGND VPWR VPWR OVHB\[6\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13750_ _13746_/CLK line[53] VGND VGND VPWR VPWR _13751_/A sky130_fd_sc_hd__dfxtp_1
X_10962_ _11032_/A VGND VGND VPWR VPWR _10962_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__05680__D line[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10298__D line[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ _12700_/Q _12712_/Y VGND VGND VPWR VPWR _13541_/Z sky130_fd_sc_hd__ebufn_2
X_10893_ _10903_/CLK line[32] VGND VGND VPWR VPWR _10893_/Q sky130_fd_sc_hd__dfxtp_1
X_13681_ _13681_/A _13692_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _12638_/CLK line[54] VGND VGND VPWR VPWR _12632_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.MUX\[14\]_A1 _05584_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12563_ _12562_/Q _12572_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13402__D line[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _11500_/CLK line[55] VGND VGND VPWR VPWR _11514_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12490_/CLK line[119] VGND VGND VPWR VPWR _12494_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11445_ _11445_/A _11452_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__09177__A _09352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[7\] clk VGND VGND VPWR VPWR _05220_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11376_ _11370_/CLK line[120] VGND VGND VPWR VPWR _11377_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10761__D line[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13115_ _13114_/Q _13132_/Y VGND VGND VPWR VPWR _11435_/Z sky130_fd_sc_hd__ebufn_2
X_10327_ _10326_/Q _10332_/Y VGND VGND VPWR VPWR _10887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05855__D line[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ _13050_/CLK line[115] VGND VGND VPWR VPWR _13046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10258_ _10248_/CLK line[121] VGND VGND VPWR VPWR _10259_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10189_ _10189_/A _10192_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[12\].TOBUF OVHB\[26\].VALID\[12\].FF/Q OVHB\[26\].INV/Y VGND VGND
+ VPWR VPWR _04933_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12688__D line[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06686__D line[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13948_ A_h[5] VGND VGND VPWR VPWR _13950_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__09062__D line[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10786__A _13932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13879_ _13879_/A _13902_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09997__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06420_ _06419_/Q _06447_/Y VGND VGND VPWR VPWR _05020_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10001__D line[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[5\] clk VGND VGND VPWR VPWR _11590_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XOVHB\[25\].VALID\[7\].FF OVHB\[25\].V/CLK A[16] VGND VGND VPWR VPWR OVHB\[25\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10936__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06351_ _06353_/CLK line[13] VGND VGND VPWR VPWR _06351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13312__D line[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05302_ _05301_/Q _05327_/Y VGND VGND VPWR VPWR _05582_/Z sky130_fd_sc_hd__ebufn_2
X_09070_ _09070_/CLK _09071_/X VGND VGND VPWR VPWR _09068_/CLK sky130_fd_sc_hd__dlclkp_1
X_06282_ _06281_/Q _06307_/Y VGND VGND VPWR VPWR _13562_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07310__D line[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08021_ _13920_/X wr VGND VGND VPWR VPWR _08021_/X sky130_fd_sc_hd__and2_1
X_05233_ _05253_/CLK line[14] VGND VGND VPWR VPWR _05233_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[4\].TOBUF OVHB\[6\].VALID\[4\].FF/Q OVHB\[6\].INV/Y VGND VGND VPWR
+ VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_7_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05164_ _05163_/Q _05187_/Y VGND VGND VPWR VPWR _05164_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09972_ _09978_/CLK line[118] VGND VGND VPWR VPWR _09973_/A sky130_fd_sc_hd__dfxtp_1
X_05095_ _05093_/CLK line[79] VGND VGND VPWR VPWR _05095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09237__D line[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08923_ _08923_/A _08932_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08854_ _08850_/CLK line[119] VGND VGND VPWR VPWR _08854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07805_ _07804_/Q _07812_/Y VGND VGND VPWR VPWR _13405_/Z sky130_fd_sc_hd__ebufn_2
X_08785_ _08784_/Q _08792_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
X_05997_ _06023_/CLK line[107] VGND VGND VPWR VPWR _05997_/Q sky130_fd_sc_hd__dfxtp_1
X_07736_ _07724_/CLK line[120] VGND VGND VPWR VPWR _07737_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06596__D line[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_04948_ _04947_/Q _04977_/Y VGND VGND VPWR VPWR _04948_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[6\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07667_ _07666_/Q _07672_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06618_ _06596_/CLK line[121] VGND VGND VPWR VPWR _06619_/A sky130_fd_sc_hd__dfxtp_1
X_09406_ _09414_/CLK line[115] VGND VGND VPWR VPWR _09406_/Q sky130_fd_sc_hd__dfxtp_1
X_07598_ _07572_/CLK line[57] VGND VGND VPWR VPWR _07598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09337_ _09336_/Q _09352_/Y VGND VGND VPWR VPWR _07097_/Z sky130_fd_sc_hd__ebufn_2
X_06549_ _06549_/A _06552_/Y VGND VGND VPWR VPWR _13549_/Z sky130_fd_sc_hd__ebufn_2
X_09268_ _09256_/CLK line[52] VGND VGND VPWR VPWR _09268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07220__D line[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08219_ _08219_/A _08232_/Y VGND VGND VPWR VPWR _06539_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09199_ _09198_/Q _09212_/Y VGND VGND VPWR VPWR _10039_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[9\].FF OVHB\[23\].V/CLK A[18] VGND VGND VPWR VPWR OVHB\[23\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11230_ _11216_/CLK line[53] VGND VGND VPWR VPWR _11230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11677__D line[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11161_ _11160_/Q _11172_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09147__D line[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10112_ _10100_/CLK line[54] VGND VGND VPWR VPWR _10112_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08051__D line[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11092_ _11090_/CLK line[118] VGND VGND VPWR VPWR _11092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13892__D line[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10043_ _10042_/Q _10052_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08986__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12151__A _12151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12301__D line[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _13822_/CLK line[91] VGND VGND VPWR VPWR _13802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11994_ _12002_/CLK line[18] VGND VGND VPWR VPWR _11994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13733_ _13733_/A _13762_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
X_10945_ _10944_/Q _10962_/Y VGND VGND VPWR VPWR _13465_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13664_ _13682_/CLK line[28] VGND VGND VPWR VPWR _13665_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09610__D line[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10876_ _10872_/CLK line[19] VGND VGND VPWR VPWR _10876_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12615_ _12614_/Q _12642_/Y VGND VGND VPWR VPWR _07015_/Z sky130_fd_sc_hd__ebufn_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13594_/Q _13622_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08226__D line[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12546_ _12560_/CLK line[29] VGND VGND VPWR VPWR _12546_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12326__A _13943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12477_ _12476_/Q _12502_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11428_ _11440_/CLK line[30] VGND VGND VPWR VPWR _11428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10491__D line[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11359_ _11358_/Q _11382_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05585__D line[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05920_ _05920_/CLK _05921_/X VGND VGND VPWR VPWR _05902_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13029_ _13028_/Q _13062_/Y VGND VGND VPWR VPWR _13589_/Z sky130_fd_sc_hd__ebufn_2
X_05851_ _13910_/X wr VGND VGND VPWR VPWR _05851_/X sky130_fd_sc_hd__and2_1
X_08570_ _08560_/CLK line[117] VGND VGND VPWR VPWR _08570_/Q sky130_fd_sc_hd__dfxtp_1
X_05782_ _13909_/X VGND VGND VPWR VPWR _05782_/Y sky130_fd_sc_hd__inv_2
X_07521_ _07520_/Q _07532_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[9\].TOBUF OVHB\[4\].VALID\[9\].FF/Q OVHB\[4\].INV/Y VGND VGND VPWR
+ VPWR _04918_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[11\].FF_D A[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[14\].VOBUF OVHB\[14\].V/Q OVHB\[14\].INV/Y VGND VGND VPWR VPWR _04916_/B1 sky130_fd_sc_hd__ebufn_2
X_07452_ _07446_/CLK line[118] VGND VGND VPWR VPWR _07452_/Q sky130_fd_sc_hd__dfxtp_1
X_06403_ _06402_/Q _06412_/Y VGND VGND VPWR VPWR _10883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10666__D line[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07383_ _07382_/Q _07392_/Y VGND VGND VPWR VPWR _06543_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13042__D line[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09122_ _09116_/CLK line[113] VGND VGND VPWR VPWR _09122_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[29\].CLKBUF\[0\]_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06334_ _06320_/CLK line[119] VGND VGND VPWR VPWR _06334_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08136__D line[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12881__D line[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09053_ _09053_/A _09072_/Y VGND VGND VPWR VPWR _06533_/Z sky130_fd_sc_hd__ebufn_2
X_06265_ _06265_/A _06272_/Y VGND VGND VPWR VPWR _06545_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07975__D line[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08004_ _08000_/CLK line[114] VGND VGND VPWR VPWR _08004_/Q sky130_fd_sc_hd__dfxtp_1
X_05216_ _05214_/CLK line[120] VGND VGND VPWR VPWR _05217_/A sky130_fd_sc_hd__dfxtp_1
X_06196_ _06186_/CLK line[56] VGND VGND VPWR VPWR _06196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05147_ _05146_/Q _05152_/Y VGND VGND VPWR VPWR _13547_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05078_ _05058_/CLK line[57] VGND VGND VPWR VPWR _05079_/A sky130_fd_sc_hd__dfxtp_1
X_09955_ _09954_/Q _09982_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08906_ _08922_/CLK line[29] VGND VGND VPWR VPWR _08907_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09886_ _09908_/CLK line[93] VGND VGND VPWR VPWR _09887_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08837_ _08837_/A _08862_/Y VGND VGND VPWR VPWR _13597_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13217__D line[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08768_ _08762_/CLK line[94] VGND VGND VPWR VPWR _08768_/Q sky130_fd_sc_hd__dfxtp_1
X_07719_ _07719_/A _07742_/Y VGND VGND VPWR VPWR _13599_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08699_ _08699_/A _08722_/Y VGND VGND VPWR VPWR _13459_/Z sky130_fd_sc_hd__ebufn_2
X_10730_ _10728_/CLK line[95] VGND VGND VPWR VPWR _10730_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].VALID\[5\].FF_D A[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10661_ _10660_/Q _10682_/Y VGND VGND VPWR VPWR _13461_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12400_ _12414_/CLK line[90] VGND VGND VPWR VPWR _12400_/Q sky130_fd_sc_hd__dfxtp_1
X_13380_ _13394_/CLK line[26] VGND VGND VPWR VPWR _13381_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10592_ _10594_/CLK line[17] VGND VGND VPWR VPWR _10592_/Q sky130_fd_sc_hd__dfxtp_1
X_12331_ _12330_/Q _12362_/Y VGND VGND VPWR VPWR _13451_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12791__D line[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[4\].TOBUF OVHB\[11\].VALID\[4\].FF/Q OVHB\[11\].INV/Y VGND VGND
+ VPWR VPWR _04939_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_103_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07885__D line[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12262_ _12268_/CLK line[27] VGND VGND VPWR VPWR _12263_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11213_ _11212_/Q _11242_/Y VGND VGND VPWR VPWR _10373_/Z sky130_fd_sc_hd__ebufn_2
X_12193_ _12193_/A _12222_/Y VGND VGND VPWR VPWR _13593_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11144_ _11148_/CLK line[28] VGND VGND VPWR VPWR _11144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11075_ _11074_/Q _11102_/Y VGND VGND VPWR VPWR _13595_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10026_ _10042_/CLK line[29] VGND VGND VPWR VPWR _10026_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12031__D line[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07125__D line[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12966__D line[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11977_ _12151_/A VGND VGND VPWR VPWR _11977_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13716_ _13715_/Q _13727_/Y VGND VGND VPWR VPWR _05036_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06964__D line[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10928_ _10930_/CLK line[48] VGND VGND VPWR VPWR _10928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09340__D line[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13647_ _13631_/CLK line[6] VGND VGND VPWR VPWR _13648_/A sky130_fd_sc_hd__dfxtp_1
X_10859_ _10858_/Q _10892_/Y VGND VGND VPWR VPWR _10859_/Z sky130_fd_sc_hd__ebufn_2
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _13577_/Q _13587_/Y VGND VGND VPWR VPWR _13578_/Z sky130_fd_sc_hd__ebufn_2
X_12529_ _12523_/CLK line[7] VGND VGND VPWR VPWR _12529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06050_ _06050_/CLK line[117] VGND VGND VPWR VPWR _06050_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[2\].FF_D A[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_MUX.MUX\[27\]_A0 _10863_/Z VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05001_ _05000_/Q _05012_/Y VGND VGND VPWR VPWR _10881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12206__D line[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09740_ _09760_/CLK line[26] VGND VGND VPWR VPWR _09740_/Q sky130_fd_sc_hd__dfxtp_1
X_06952_ _06960_/CLK line[17] VGND VGND VPWR VPWR _06952_/Q sky130_fd_sc_hd__dfxtp_1
.ends

