VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM
  CLASS BLOCK ;
  FOREIGN DFFRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 1089.200 BY 1389.360 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.460 1385.360 452.740 1389.360 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.720 1385.360 467.000 1389.360 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.980 1385.360 481.260 1389.360 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.780 1385.360 495.060 1389.360 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.040 1385.360 509.320 1389.360 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.300 1385.360 523.580 1389.360 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.100 1385.360 537.380 1389.360 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.360 1385.360 551.640 1389.360 ;
    END
  END A[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.620 1385.360 565.900 1389.360 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.260 1385.360 650.540 1389.360 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.020 1385.360 791.300 1389.360 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.280 1385.360 805.560 1389.360 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.080 1385.360 819.360 1389.360 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.340 1385.360 833.620 1389.360 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.600 1385.360 847.880 1389.360 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.400 1385.360 861.680 1389.360 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.660 1385.360 875.940 1389.360 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.920 1385.360 890.200 1389.360 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.720 1385.360 904.000 1389.360 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.980 1385.360 918.260 1389.360 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.060 1385.360 664.340 1389.360 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.240 1385.360 932.520 1389.360 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.040 1385.360 946.320 1389.360 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.300 1385.360 960.580 1389.360 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.560 1385.360 974.840 1389.360 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.360 1385.360 988.640 1389.360 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.620 1385.360 1002.900 1389.360 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.880 1385.360 1017.160 1389.360 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.680 1385.360 1030.960 1389.360 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.940 1385.360 1045.220 1389.360 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.200 1385.360 1059.480 1389.360 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.320 1385.360 678.600 1389.360 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.000 1385.360 1073.280 1389.360 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.260 1385.360 1087.540 1389.360 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.580 1385.360 692.860 1389.360 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.380 1385.360 706.660 1389.360 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.640 1385.360 720.920 1389.360 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.900 1385.360 735.180 1389.360 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.700 1385.360 748.980 1389.360 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.960 1385.360 763.240 1389.360 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.760 1385.360 777.040 1389.360 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.660 1385.360 1.940 1389.360 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.420 1385.360 142.700 1389.360 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.680 1385.360 156.960 1389.360 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.480 1385.360 170.760 1389.360 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.740 1385.360 185.020 1389.360 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.000 1385.360 199.280 1389.360 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.800 1385.360 213.080 1389.360 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.060 1385.360 227.340 1389.360 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.320 1385.360 241.600 1389.360 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.120 1385.360 255.400 1389.360 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.380 1385.360 269.660 1389.360 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.460 1385.360 15.740 1389.360 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.640 1385.360 283.920 1389.360 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.440 1385.360 297.720 1389.360 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.700 1385.360 311.980 1389.360 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.960 1385.360 326.240 1389.360 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.760 1385.360 340.040 1389.360 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.020 1385.360 354.300 1389.360 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.280 1385.360 368.560 1389.360 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.080 1385.360 382.360 1389.360 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.340 1385.360 396.620 1389.360 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.140 1385.360 410.420 1389.360 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.720 1385.360 30.000 1389.360 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.400 1385.360 424.680 1389.360 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.660 1385.360 438.940 1389.360 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.520 1385.360 43.800 1389.360 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.780 1385.360 58.060 1389.360 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.040 1385.360 72.320 1389.360 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.840 1385.360 86.120 1389.360 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.100 1385.360 100.380 1389.360 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.360 1385.360 114.640 1389.360 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.160 1385.360 128.440 1389.360 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.000 1385.360 636.280 1389.360 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.420 1385.360 579.700 1389.360 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.680 1385.360 593.960 1389.360 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.940 1385.360 608.220 1389.360 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.740 1385.360 622.020 1389.360 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.310 0.000 938.910 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.710 0.000 785.310 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 630.110 0.000 631.710 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 476.510 0.000 478.110 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 322.910 0.000 324.510 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 169.310 0.000 170.910 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 0.000 17.310 1376.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1014.110 0.000 1015.710 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 860.510 0.000 862.110 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.910 0.000 708.510 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 553.310 0.000 554.910 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 399.710 0.000 401.310 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.110 0.000 247.710 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 0.000 94.110 1376.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 0.155 1089.010 1376.645 ;
      LAYER met1 ;
        RECT 0.190 0.000 1089.010 1377.200 ;
      LAYER met2 ;
        RECT 2.220 1385.080 15.180 1385.360 ;
        RECT 16.020 1385.080 29.440 1385.360 ;
        RECT 30.280 1385.080 43.240 1385.360 ;
        RECT 44.080 1385.080 57.500 1385.360 ;
        RECT 58.340 1385.080 71.760 1385.360 ;
        RECT 72.600 1385.080 85.560 1385.360 ;
        RECT 86.400 1385.080 99.820 1385.360 ;
        RECT 100.660 1385.080 114.080 1385.360 ;
        RECT 114.920 1385.080 127.880 1385.360 ;
        RECT 128.720 1385.080 142.140 1385.360 ;
        RECT 142.980 1385.080 156.400 1385.360 ;
        RECT 157.240 1385.080 170.200 1385.360 ;
        RECT 171.040 1385.080 184.460 1385.360 ;
        RECT 185.300 1385.080 198.720 1385.360 ;
        RECT 199.560 1385.080 212.520 1385.360 ;
        RECT 213.360 1385.080 226.780 1385.360 ;
        RECT 227.620 1385.080 241.040 1385.360 ;
        RECT 241.880 1385.080 254.840 1385.360 ;
        RECT 255.680 1385.080 269.100 1385.360 ;
        RECT 269.940 1385.080 283.360 1385.360 ;
        RECT 284.200 1385.080 297.160 1385.360 ;
        RECT 298.000 1385.080 311.420 1385.360 ;
        RECT 312.260 1385.080 325.680 1385.360 ;
        RECT 326.520 1385.080 339.480 1385.360 ;
        RECT 340.320 1385.080 353.740 1385.360 ;
        RECT 354.580 1385.080 368.000 1385.360 ;
        RECT 368.840 1385.080 381.800 1385.360 ;
        RECT 382.640 1385.080 396.060 1385.360 ;
        RECT 396.900 1385.080 409.860 1385.360 ;
        RECT 410.700 1385.080 424.120 1385.360 ;
        RECT 424.960 1385.080 438.380 1385.360 ;
        RECT 439.220 1385.080 452.180 1385.360 ;
        RECT 453.020 1385.080 466.440 1385.360 ;
        RECT 467.280 1385.080 480.700 1385.360 ;
        RECT 481.540 1385.080 494.500 1385.360 ;
        RECT 495.340 1385.080 508.760 1385.360 ;
        RECT 509.600 1385.080 523.020 1385.360 ;
        RECT 523.860 1385.080 536.820 1385.360 ;
        RECT 537.660 1385.080 551.080 1385.360 ;
        RECT 551.920 1385.080 565.340 1385.360 ;
        RECT 566.180 1385.080 579.140 1385.360 ;
        RECT 579.980 1385.080 593.400 1385.360 ;
        RECT 594.240 1385.080 607.660 1385.360 ;
        RECT 608.500 1385.080 621.460 1385.360 ;
        RECT 622.300 1385.080 635.720 1385.360 ;
        RECT 636.560 1385.080 649.980 1385.360 ;
        RECT 650.820 1385.080 663.780 1385.360 ;
        RECT 664.620 1385.080 678.040 1385.360 ;
        RECT 678.880 1385.080 692.300 1385.360 ;
        RECT 693.140 1385.080 706.100 1385.360 ;
        RECT 706.940 1385.080 720.360 1385.360 ;
        RECT 721.200 1385.080 734.620 1385.360 ;
        RECT 735.460 1385.080 748.420 1385.360 ;
        RECT 749.260 1385.080 762.680 1385.360 ;
        RECT 763.520 1385.080 776.480 1385.360 ;
        RECT 777.320 1385.080 790.740 1385.360 ;
        RECT 791.580 1385.080 805.000 1385.360 ;
        RECT 805.840 1385.080 818.800 1385.360 ;
        RECT 819.640 1385.080 833.060 1385.360 ;
        RECT 833.900 1385.080 847.320 1385.360 ;
        RECT 848.160 1385.080 861.120 1385.360 ;
        RECT 861.960 1385.080 875.380 1385.360 ;
        RECT 876.220 1385.080 889.640 1385.360 ;
        RECT 890.480 1385.080 903.440 1385.360 ;
        RECT 904.280 1385.080 917.700 1385.360 ;
        RECT 918.540 1385.080 931.960 1385.360 ;
        RECT 932.800 1385.080 945.760 1385.360 ;
        RECT 946.600 1385.080 960.020 1385.360 ;
        RECT 960.860 1385.080 974.280 1385.360 ;
        RECT 975.120 1385.080 988.080 1385.360 ;
        RECT 988.920 1385.080 1002.340 1385.360 ;
        RECT 1003.180 1385.080 1016.600 1385.360 ;
        RECT 1017.440 1385.080 1030.400 1385.360 ;
        RECT 1031.240 1385.080 1044.660 1385.360 ;
        RECT 1045.500 1385.080 1058.920 1385.360 ;
        RECT 1059.760 1385.080 1072.720 1385.360 ;
        RECT 1073.560 1385.080 1086.980 1385.360 ;
        RECT 1.670 0.000 1087.530 1385.080 ;
      LAYER met3 ;
        RECT 4.395 0.075 1015.710 1376.725 ;
      LAYER met4 ;
        RECT 139.405 753.175 168.910 1374.345 ;
        RECT 171.310 753.175 245.710 1374.345 ;
        RECT 248.110 753.175 322.510 1374.345 ;
        RECT 324.910 753.175 399.310 1374.345 ;
        RECT 401.710 753.175 476.110 1374.345 ;
        RECT 478.510 753.175 552.910 1374.345 ;
        RECT 555.310 753.175 629.710 1374.345 ;
        RECT 632.110 753.175 706.510 1374.345 ;
        RECT 708.910 753.175 783.310 1374.345 ;
        RECT 785.710 753.175 846.295 1374.345 ;
  END
END DFFRAM
END LIBRARY

