magic
tech sky130A
magscale 1 2
timestamp 1609364000
<< obsli1 >>
rect 38 31 217957 275329
<< obsm1 >>
rect 38 0 217969 276052
<< metal2 >>
rect 240 277072 296 277872
rect 2908 277072 2964 277872
rect 5668 277072 5724 277872
rect 8428 277072 8484 277872
rect 11188 277072 11244 277872
rect 13948 277072 14004 277872
rect 16708 277072 16764 277872
rect 19468 277072 19524 277872
rect 22228 277072 22284 277872
rect 24896 277072 24952 277872
rect 27656 277072 27712 277872
rect 30416 277072 30472 277872
rect 33176 277072 33232 277872
rect 35936 277072 35992 277872
rect 38696 277072 38752 277872
rect 41456 277072 41512 277872
rect 44216 277072 44272 277872
rect 46976 277072 47032 277872
rect 49644 277072 49700 277872
rect 52404 277072 52460 277872
rect 55164 277072 55220 277872
rect 57924 277072 57980 277872
rect 60684 277072 60740 277872
rect 63444 277072 63500 277872
rect 66204 277072 66260 277872
rect 68964 277072 69020 277872
rect 71724 277072 71780 277872
rect 74392 277072 74448 277872
rect 77152 277072 77208 277872
rect 79912 277072 79968 277872
rect 82672 277072 82728 277872
rect 85432 277072 85488 277872
rect 88192 277072 88248 277872
rect 90952 277072 91008 277872
rect 93712 277072 93768 277872
rect 96472 277072 96528 277872
rect 99140 277072 99196 277872
rect 101900 277072 101956 277872
rect 104660 277072 104716 277872
rect 107420 277072 107476 277872
rect 110180 277072 110236 277872
rect 112940 277072 112996 277872
rect 115700 277072 115756 277872
rect 118460 277072 118516 277872
rect 121220 277072 121276 277872
rect 123888 277072 123944 277872
rect 126648 277072 126704 277872
rect 129408 277072 129464 277872
rect 132168 277072 132224 277872
rect 134928 277072 134984 277872
rect 137688 277072 137744 277872
rect 140448 277072 140504 277872
rect 143208 277072 143264 277872
rect 145968 277072 146024 277872
rect 148636 277072 148692 277872
rect 151396 277072 151452 277872
rect 154156 277072 154212 277872
rect 156916 277072 156972 277872
rect 159676 277072 159732 277872
rect 162436 277072 162492 277872
rect 165196 277072 165252 277872
rect 167956 277072 168012 277872
rect 170716 277072 170772 277872
rect 173384 277072 173440 277872
rect 176144 277072 176200 277872
rect 178904 277072 178960 277872
rect 181664 277072 181720 277872
rect 184424 277072 184480 277872
rect 187184 277072 187240 277872
rect 189944 277072 190000 277872
rect 192704 277072 192760 277872
rect 195464 277072 195520 277872
rect 198132 277072 198188 277872
rect 200892 277072 200948 277872
rect 203652 277072 203708 277872
rect 206412 277072 206468 277872
rect 209172 277072 209228 277872
rect 211932 277072 211988 277872
rect 214692 277072 214748 277872
rect 217452 277072 217508 277872
<< obsm2 >>
rect 352 277016 2852 277072
rect 3020 277016 5612 277072
rect 5780 277016 8372 277072
rect 8540 277016 11132 277072
rect 11300 277016 13892 277072
rect 14060 277016 16652 277072
rect 16820 277016 19412 277072
rect 19580 277016 22172 277072
rect 22340 277016 24840 277072
rect 25008 277016 27600 277072
rect 27768 277016 30360 277072
rect 30528 277016 33120 277072
rect 33288 277016 35880 277072
rect 36048 277016 38640 277072
rect 38808 277016 41400 277072
rect 41568 277016 44160 277072
rect 44328 277016 46920 277072
rect 47088 277016 49588 277072
rect 49756 277016 52348 277072
rect 52516 277016 55108 277072
rect 55276 277016 57868 277072
rect 58036 277016 60628 277072
rect 60796 277016 63388 277072
rect 63556 277016 66148 277072
rect 66316 277016 68908 277072
rect 69076 277016 71668 277072
rect 71836 277016 74336 277072
rect 74504 277016 77096 277072
rect 77264 277016 79856 277072
rect 80024 277016 82616 277072
rect 82784 277016 85376 277072
rect 85544 277016 88136 277072
rect 88304 277016 90896 277072
rect 91064 277016 93656 277072
rect 93824 277016 96416 277072
rect 96584 277016 99084 277072
rect 99252 277016 101844 277072
rect 102012 277016 104604 277072
rect 104772 277016 107364 277072
rect 107532 277016 110124 277072
rect 110292 277016 112884 277072
rect 113052 277016 115644 277072
rect 115812 277016 118404 277072
rect 118572 277016 121164 277072
rect 121332 277016 123832 277072
rect 124000 277016 126592 277072
rect 126760 277016 129352 277072
rect 129520 277016 132112 277072
rect 132280 277016 134872 277072
rect 135040 277016 137632 277072
rect 137800 277016 140392 277072
rect 140560 277016 143152 277072
rect 143320 277016 145912 277072
rect 146080 277016 148580 277072
rect 148748 277016 151340 277072
rect 151508 277016 154100 277072
rect 154268 277016 156860 277072
rect 157028 277016 159620 277072
rect 159788 277016 162380 277072
rect 162548 277016 165140 277072
rect 165308 277016 167900 277072
rect 168068 277016 170660 277072
rect 170828 277016 173328 277072
rect 173496 277016 176088 277072
rect 176256 277016 178848 277072
rect 179016 277016 181608 277072
rect 181776 277016 184368 277072
rect 184536 277016 187128 277072
rect 187296 277016 189888 277072
rect 190056 277016 192648 277072
rect 192816 277016 195408 277072
rect 195576 277016 198076 277072
rect 198244 277016 200836 277072
rect 201004 277016 203596 277072
rect 203764 277016 206356 277072
rect 206524 277016 209116 277072
rect 209284 277016 211876 277072
rect 212044 277016 214636 277072
rect 214804 277016 217396 277072
rect 217564 277016 217600 277072
rect 242 0 217600 277016
<< obsm3 >>
rect 327 15 217605 275345
<< metal4 >>
rect 3142 0 3462 275360
rect 18502 0 18822 275360
rect 33862 0 34182 275360
rect 49222 0 49542 275360
rect 64582 0 64902 275360
rect 79942 0 80262 275360
rect 95302 0 95622 275360
rect 110662 0 110982 275360
rect 126022 0 126342 275360
rect 141382 0 141702 275360
rect 156742 0 157062 275360
rect 172102 0 172422 275360
rect 187462 0 187782 275360
rect 202822 0 203142 275360
<< obsm4 >>
rect 2305 3891 3062 275005
rect 3542 3891 18422 275005
rect 18902 3891 33782 275005
rect 34262 3891 49142 275005
rect 49622 3891 64502 275005
rect 64982 3891 79862 275005
rect 80342 3891 95222 275005
rect 95702 3891 110582 275005
rect 111062 3891 125942 275005
rect 126422 3891 141302 275005
rect 141782 3891 156662 275005
rect 157142 3891 172022 275005
rect 172502 3891 187382 275005
rect 187862 3891 202742 275005
rect 203222 3891 213971 275005
<< labels >>
rlabel metal2 s 88192 277072 88248 277872 6 A[0]
port 1 nsew signal input
rlabel metal2 s 90952 277072 91008 277872 6 A[1]
port 2 nsew signal input
rlabel metal2 s 93712 277072 93768 277872 6 A[2]
port 3 nsew signal input
rlabel metal2 s 96472 277072 96528 277872 6 A[3]
port 4 nsew signal input
rlabel metal2 s 99140 277072 99196 277872 6 A[4]
port 5 nsew signal input
rlabel metal2 s 101900 277072 101956 277872 6 A[5]
port 6 nsew signal input
rlabel metal2 s 104660 277072 104716 277872 6 A[6]
port 7 nsew signal input
rlabel metal2 s 107420 277072 107476 277872 6 A[7]
port 8 nsew signal input
rlabel metal2 s 110180 277072 110236 277872 6 A[8]
port 9 nsew signal input
rlabel metal2 s 112940 277072 112996 277872 6 A[9]
port 10 nsew signal input
rlabel metal2 s 115700 277072 115756 277872 6 CLK
port 11 nsew signal input
rlabel metal2 s 132168 277072 132224 277872 6 Di[0]
port 12 nsew signal input
rlabel metal2 s 159676 277072 159732 277872 6 Di[10]
port 13 nsew signal input
rlabel metal2 s 162436 277072 162492 277872 6 Di[11]
port 14 nsew signal input
rlabel metal2 s 165196 277072 165252 277872 6 Di[12]
port 15 nsew signal input
rlabel metal2 s 167956 277072 168012 277872 6 Di[13]
port 16 nsew signal input
rlabel metal2 s 170716 277072 170772 277872 6 Di[14]
port 17 nsew signal input
rlabel metal2 s 173384 277072 173440 277872 6 Di[15]
port 18 nsew signal input
rlabel metal2 s 176144 277072 176200 277872 6 Di[16]
port 19 nsew signal input
rlabel metal2 s 178904 277072 178960 277872 6 Di[17]
port 20 nsew signal input
rlabel metal2 s 181664 277072 181720 277872 6 Di[18]
port 21 nsew signal input
rlabel metal2 s 184424 277072 184480 277872 6 Di[19]
port 22 nsew signal input
rlabel metal2 s 134928 277072 134984 277872 6 Di[1]
port 23 nsew signal input
rlabel metal2 s 187184 277072 187240 277872 6 Di[20]
port 24 nsew signal input
rlabel metal2 s 189944 277072 190000 277872 6 Di[21]
port 25 nsew signal input
rlabel metal2 s 192704 277072 192760 277872 6 Di[22]
port 26 nsew signal input
rlabel metal2 s 195464 277072 195520 277872 6 Di[23]
port 27 nsew signal input
rlabel metal2 s 198132 277072 198188 277872 6 Di[24]
port 28 nsew signal input
rlabel metal2 s 200892 277072 200948 277872 6 Di[25]
port 29 nsew signal input
rlabel metal2 s 203652 277072 203708 277872 6 Di[26]
port 30 nsew signal input
rlabel metal2 s 206412 277072 206468 277872 6 Di[27]
port 31 nsew signal input
rlabel metal2 s 209172 277072 209228 277872 6 Di[28]
port 32 nsew signal input
rlabel metal2 s 211932 277072 211988 277872 6 Di[29]
port 33 nsew signal input
rlabel metal2 s 137688 277072 137744 277872 6 Di[2]
port 34 nsew signal input
rlabel metal2 s 214692 277072 214748 277872 6 Di[30]
port 35 nsew signal input
rlabel metal2 s 217452 277072 217508 277872 6 Di[31]
port 36 nsew signal input
rlabel metal2 s 140448 277072 140504 277872 6 Di[3]
port 37 nsew signal input
rlabel metal2 s 143208 277072 143264 277872 6 Di[4]
port 38 nsew signal input
rlabel metal2 s 145968 277072 146024 277872 6 Di[5]
port 39 nsew signal input
rlabel metal2 s 148636 277072 148692 277872 6 Di[6]
port 40 nsew signal input
rlabel metal2 s 151396 277072 151452 277872 6 Di[7]
port 41 nsew signal input
rlabel metal2 s 154156 277072 154212 277872 6 Di[8]
port 42 nsew signal input
rlabel metal2 s 156916 277072 156972 277872 6 Di[9]
port 43 nsew signal input
rlabel metal2 s 240 277072 296 277872 6 Do[0]
port 44 nsew signal output
rlabel metal2 s 27656 277072 27712 277872 6 Do[10]
port 45 nsew signal output
rlabel metal2 s 30416 277072 30472 277872 6 Do[11]
port 46 nsew signal output
rlabel metal2 s 33176 277072 33232 277872 6 Do[12]
port 47 nsew signal output
rlabel metal2 s 35936 277072 35992 277872 6 Do[13]
port 48 nsew signal output
rlabel metal2 s 38696 277072 38752 277872 6 Do[14]
port 49 nsew signal output
rlabel metal2 s 41456 277072 41512 277872 6 Do[15]
port 50 nsew signal output
rlabel metal2 s 44216 277072 44272 277872 6 Do[16]
port 51 nsew signal output
rlabel metal2 s 46976 277072 47032 277872 6 Do[17]
port 52 nsew signal output
rlabel metal2 s 49644 277072 49700 277872 6 Do[18]
port 53 nsew signal output
rlabel metal2 s 52404 277072 52460 277872 6 Do[19]
port 54 nsew signal output
rlabel metal2 s 2908 277072 2964 277872 6 Do[1]
port 55 nsew signal output
rlabel metal2 s 55164 277072 55220 277872 6 Do[20]
port 56 nsew signal output
rlabel metal2 s 57924 277072 57980 277872 6 Do[21]
port 57 nsew signal output
rlabel metal2 s 60684 277072 60740 277872 6 Do[22]
port 58 nsew signal output
rlabel metal2 s 63444 277072 63500 277872 6 Do[23]
port 59 nsew signal output
rlabel metal2 s 66204 277072 66260 277872 6 Do[24]
port 60 nsew signal output
rlabel metal2 s 68964 277072 69020 277872 6 Do[25]
port 61 nsew signal output
rlabel metal2 s 71724 277072 71780 277872 6 Do[26]
port 62 nsew signal output
rlabel metal2 s 74392 277072 74448 277872 6 Do[27]
port 63 nsew signal output
rlabel metal2 s 77152 277072 77208 277872 6 Do[28]
port 64 nsew signal output
rlabel metal2 s 79912 277072 79968 277872 6 Do[29]
port 65 nsew signal output
rlabel metal2 s 5668 277072 5724 277872 6 Do[2]
port 66 nsew signal output
rlabel metal2 s 82672 277072 82728 277872 6 Do[30]
port 67 nsew signal output
rlabel metal2 s 85432 277072 85488 277872 6 Do[31]
port 68 nsew signal output
rlabel metal2 s 8428 277072 8484 277872 6 Do[3]
port 69 nsew signal output
rlabel metal2 s 11188 277072 11244 277872 6 Do[4]
port 70 nsew signal output
rlabel metal2 s 13948 277072 14004 277872 6 Do[5]
port 71 nsew signal output
rlabel metal2 s 16708 277072 16764 277872 6 Do[6]
port 72 nsew signal output
rlabel metal2 s 19468 277072 19524 277872 6 Do[7]
port 73 nsew signal output
rlabel metal2 s 22228 277072 22284 277872 6 Do[8]
port 74 nsew signal output
rlabel metal2 s 24896 277072 24952 277872 6 Do[9]
port 75 nsew signal output
rlabel metal2 s 129408 277072 129464 277872 6 EN
port 76 nsew signal input
rlabel metal2 s 118460 277072 118516 277872 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 121220 277072 121276 277872 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 123888 277072 123944 277872 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 126648 277072 126704 277872 6 WE[3]
port 80 nsew signal input
rlabel metal4 s 187462 0 187782 275360 6 VPWR
port 81 nsew power bidirectional
rlabel metal4 s 156742 0 157062 275360 6 VPWR
port 82 nsew power bidirectional
rlabel metal4 s 126022 0 126342 275360 6 VPWR
port 83 nsew power bidirectional
rlabel metal4 s 95302 0 95622 275360 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 64582 0 64902 275360 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 33862 0 34182 275360 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 3142 0 3462 275360 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 202822 0 203142 275360 6 VGND
port 88 nsew ground bidirectional
rlabel metal4 s 172102 0 172422 275360 6 VGND
port 89 nsew ground bidirectional
rlabel metal4 s 141382 0 141702 275360 6 VGND
port 90 nsew ground bidirectional
rlabel metal4 s 110662 0 110982 275360 6 VGND
port 91 nsew ground bidirectional
rlabel metal4 s 79942 0 80262 275360 6 VGND
port 92 nsew ground bidirectional
rlabel metal4 s 49222 0 49542 275360 6 VGND
port 93 nsew ground bidirectional
rlabel metal4 s 18502 0 18822 275360 6 VGND
port 94 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 217969 277872
string LEFview TRUE
<< end >>
