magic
tech sky130A
magscale 1 2
timestamp 1608998679
<< obsli1 >>
rect 626 2159 78521 117521
<< obsm1 >>
rect 626 1232 78628 119128
<< metal2 >>
rect 0 119200 56 120000
rect 920 119200 976 120000
rect 1932 119200 1988 120000
rect 2944 119200 3000 120000
rect 3956 119200 4012 120000
rect 4968 119200 5024 120000
rect 5980 119200 6036 120000
rect 6992 119200 7048 120000
rect 8004 119200 8060 120000
rect 8924 119200 8980 120000
rect 9936 119200 9992 120000
rect 10948 119200 11004 120000
rect 11960 119200 12016 120000
rect 12972 119200 13028 120000
rect 13984 119200 14040 120000
rect 14996 119200 15052 120000
rect 16008 119200 16064 120000
rect 16928 119200 16984 120000
rect 17940 119200 17996 120000
rect 18952 119200 19008 120000
rect 19964 119200 20020 120000
rect 20976 119200 21032 120000
rect 21988 119200 22044 120000
rect 23000 119200 23056 120000
rect 24012 119200 24068 120000
rect 24932 119200 24988 120000
rect 25944 119200 26000 120000
rect 26956 119200 27012 120000
rect 27968 119200 28024 120000
rect 28980 119200 29036 120000
rect 29992 119200 30048 120000
rect 31004 119200 31060 120000
rect 32016 119200 32072 120000
rect 32936 119200 32992 120000
rect 33948 119200 34004 120000
rect 34960 119200 35016 120000
rect 35972 119200 36028 120000
rect 36984 119200 37040 120000
rect 37996 119200 38052 120000
rect 39008 119200 39064 120000
rect 40020 119200 40076 120000
rect 40940 119200 40996 120000
rect 41952 119200 42008 120000
rect 42964 119200 43020 120000
rect 43976 119200 44032 120000
rect 44988 119200 45044 120000
rect 46000 119200 46056 120000
rect 47012 119200 47068 120000
rect 48024 119200 48080 120000
rect 48944 119200 49000 120000
rect 49956 119200 50012 120000
rect 50968 119200 51024 120000
rect 51980 119200 52036 120000
rect 52992 119200 53048 120000
rect 54004 119200 54060 120000
rect 55016 119200 55072 120000
rect 56028 119200 56084 120000
rect 56948 119200 57004 120000
rect 57960 119200 58016 120000
rect 58972 119200 59028 120000
rect 59984 119200 60040 120000
rect 60996 119200 61052 120000
rect 62008 119200 62064 120000
rect 63020 119200 63076 120000
rect 64032 119200 64088 120000
rect 64952 119200 65008 120000
rect 65964 119200 66020 120000
rect 66976 119200 67032 120000
rect 67988 119200 68044 120000
rect 69000 119200 69056 120000
rect 70012 119200 70068 120000
rect 71024 119200 71080 120000
rect 72036 119200 72092 120000
rect 72956 119200 73012 120000
rect 73968 119200 74024 120000
rect 74980 119200 75036 120000
rect 75992 119200 76048 120000
rect 77004 119200 77060 120000
rect 78016 119200 78072 120000
rect 79028 119200 79084 120000
rect 9476 0 9532 800
rect 29440 0 29496 800
rect 49496 0 49552 800
rect 69460 0 69516 800
<< obsm2 >>
rect 1032 119144 1876 119513
rect 2044 119144 2888 119513
rect 3056 119144 3900 119513
rect 4068 119144 4912 119513
rect 5080 119144 5924 119513
rect 6092 119144 6936 119513
rect 7104 119144 7948 119513
rect 8116 119144 8868 119513
rect 9036 119144 9880 119513
rect 10048 119144 10892 119513
rect 11060 119144 11904 119513
rect 12072 119144 12916 119513
rect 13084 119144 13928 119513
rect 14096 119144 14940 119513
rect 15108 119144 15952 119513
rect 16120 119144 16872 119513
rect 17040 119144 17884 119513
rect 18052 119144 18896 119513
rect 19064 119144 19908 119513
rect 20076 119144 20920 119513
rect 21088 119144 21932 119513
rect 22100 119144 22944 119513
rect 23112 119144 23956 119513
rect 24124 119144 24876 119513
rect 25044 119144 25888 119513
rect 26056 119144 26900 119513
rect 27068 119144 27912 119513
rect 28080 119144 28924 119513
rect 29092 119144 29936 119513
rect 30104 119144 30948 119513
rect 31116 119144 31960 119513
rect 32128 119144 32880 119513
rect 33048 119144 33892 119513
rect 34060 119144 34904 119513
rect 35072 119144 35916 119513
rect 36084 119144 36928 119513
rect 37096 119144 37940 119513
rect 38108 119144 38952 119513
rect 39120 119144 39964 119513
rect 40132 119144 40884 119513
rect 41052 119144 41896 119513
rect 42064 119144 42908 119513
rect 43076 119144 43920 119513
rect 44088 119144 44932 119513
rect 45100 119144 45944 119513
rect 46112 119144 46956 119513
rect 47124 119144 47968 119513
rect 48136 119144 48888 119513
rect 49056 119144 49900 119513
rect 50068 119144 50912 119513
rect 51080 119144 51924 119513
rect 52092 119144 52936 119513
rect 53104 119144 53948 119513
rect 54116 119144 54960 119513
rect 55128 119144 55972 119513
rect 56140 119144 56892 119513
rect 57060 119144 57904 119513
rect 58072 119144 58916 119513
rect 59084 119144 59928 119513
rect 60096 119144 60940 119513
rect 61108 119144 61952 119513
rect 62120 119144 62964 119513
rect 63132 119144 63976 119513
rect 64144 119144 64896 119513
rect 65064 119144 65908 119513
rect 66076 119144 66920 119513
rect 67088 119144 67932 119513
rect 68100 119144 68944 119513
rect 69112 119144 69956 119513
rect 70124 119144 70968 119513
rect 71136 119144 71980 119513
rect 72148 119144 72900 119513
rect 73068 119144 73912 119513
rect 74080 119144 74924 119513
rect 75092 119144 75936 119513
rect 76104 119144 76948 119513
rect 77116 119144 77960 119513
rect 78128 119144 78972 119513
rect 920 856 79070 119144
rect 920 439 9420 856
rect 9588 439 29384 856
rect 29552 439 49440 856
rect 49608 439 69404 856
rect 69572 439 79070 856
<< metal3 >>
rect 78722 119416 79522 119536
rect 78722 118464 79522 118584
rect 78722 117512 79522 117632
rect 78722 116560 79522 116680
rect 78722 115608 79522 115728
rect 78722 114656 79522 114776
rect 78722 113704 79522 113824
rect 78722 112752 79522 112872
rect 78722 111800 79522 111920
rect 78722 110984 79522 111104
rect 78722 110032 79522 110152
rect 78722 109080 79522 109200
rect 78722 108128 79522 108248
rect 78722 107176 79522 107296
rect 78722 106224 79522 106344
rect 78722 105272 79522 105392
rect 78722 104320 79522 104440
rect 78722 103368 79522 103488
rect 78722 102552 79522 102672
rect 78722 101600 79522 101720
rect 78722 100648 79522 100768
rect 78722 99696 79522 99816
rect 78722 98744 79522 98864
rect 78722 97792 79522 97912
rect 78722 96840 79522 96960
rect 78722 95888 79522 96008
rect 78722 94936 79522 95056
rect 78722 94120 79522 94240
rect 78722 93168 79522 93288
rect 78722 92216 79522 92336
rect 78722 91264 79522 91384
rect 78722 90312 79522 90432
rect 78722 89360 79522 89480
rect 78722 88408 79522 88528
rect 78722 87456 79522 87576
rect 78722 86504 79522 86624
rect 78722 85688 79522 85808
rect 78722 84736 79522 84856
rect 78722 83784 79522 83904
rect 78722 82832 79522 82952
rect 78722 81880 79522 82000
rect 78722 80928 79522 81048
rect 78722 79976 79522 80096
rect 78722 79024 79522 79144
rect 78722 78072 79522 78192
rect 78722 77256 79522 77376
rect 78722 76304 79522 76424
rect 78722 75352 79522 75472
rect 78722 74400 79522 74520
rect 78722 73448 79522 73568
rect 78722 72496 79522 72616
rect 78722 71544 79522 71664
rect 78722 70592 79522 70712
rect 78722 69640 79522 69760
rect 78722 68824 79522 68944
rect 78722 67872 79522 67992
rect 78722 66920 79522 67040
rect 78722 65968 79522 66088
rect 78722 65016 79522 65136
rect 78722 64064 79522 64184
rect 78722 63112 79522 63232
rect 78722 62160 79522 62280
rect 78722 61208 79522 61328
rect 78722 60392 79522 60512
rect 78722 59440 79522 59560
rect 78722 58488 79522 58608
rect 78722 57536 79522 57656
rect 78722 56584 79522 56704
rect 78722 55632 79522 55752
rect 78722 54680 79522 54800
rect 78722 53728 79522 53848
rect 78722 52776 79522 52896
rect 78722 51824 79522 51944
rect 78722 51008 79522 51128
rect 78722 50056 79522 50176
rect 78722 49104 79522 49224
rect 78722 48152 79522 48272
rect 78722 47200 79522 47320
rect 78722 46248 79522 46368
rect 78722 45296 79522 45416
rect 78722 44344 79522 44464
rect 78722 43392 79522 43512
rect 78722 42576 79522 42696
rect 78722 41624 79522 41744
rect 78722 40672 79522 40792
rect 78722 39720 79522 39840
rect 78722 38768 79522 38888
rect 78722 37816 79522 37936
rect 78722 36864 79522 36984
rect 78722 35912 79522 36032
rect 78722 34960 79522 35080
rect 78722 34144 79522 34264
rect 78722 33192 79522 33312
rect 78722 32240 79522 32360
rect 78722 31288 79522 31408
rect 78722 30336 79522 30456
rect 78722 29384 79522 29504
rect 78722 28432 79522 28552
rect 78722 27480 79522 27600
rect 78722 26528 79522 26648
rect 78722 25712 79522 25832
rect 78722 24760 79522 24880
rect 78722 23808 79522 23928
rect 78722 22856 79522 22976
rect 78722 21904 79522 22024
rect 78722 20952 79522 21072
rect 78722 20000 79522 20120
rect 78722 19048 79522 19168
rect 78722 18096 79522 18216
rect 78722 17280 79522 17400
rect 78722 16328 79522 16448
rect 78722 15376 79522 15496
rect 78722 14424 79522 14544
rect 78722 13472 79522 13592
rect 78722 12520 79522 12640
rect 78722 11568 79522 11688
rect 78722 10616 79522 10736
rect 78722 9664 79522 9784
rect 78722 8848 79522 8968
rect 78722 7896 79522 8016
rect 78722 6944 79522 7064
rect 78722 5992 79522 6112
rect 78722 5040 79522 5160
rect 78722 4088 79522 4208
rect 78722 3136 79522 3256
rect 78722 2184 79522 2304
rect 78722 1232 79522 1352
rect 78722 416 79522 536
<< obsm3 >>
rect 915 119336 78642 119509
rect 915 118664 78722 119336
rect 915 118384 78642 118664
rect 915 117712 78722 118384
rect 915 117432 78642 117712
rect 915 116760 78722 117432
rect 915 116480 78642 116760
rect 915 115808 78722 116480
rect 915 115528 78642 115808
rect 915 114856 78722 115528
rect 915 114576 78642 114856
rect 915 113904 78722 114576
rect 915 113624 78642 113904
rect 915 112952 78722 113624
rect 915 112672 78642 112952
rect 915 112000 78722 112672
rect 915 111720 78642 112000
rect 915 111184 78722 111720
rect 915 110904 78642 111184
rect 915 110232 78722 110904
rect 915 109952 78642 110232
rect 915 109280 78722 109952
rect 915 109000 78642 109280
rect 915 108328 78722 109000
rect 915 108048 78642 108328
rect 915 107376 78722 108048
rect 915 107096 78642 107376
rect 915 106424 78722 107096
rect 915 106144 78642 106424
rect 915 105472 78722 106144
rect 915 105192 78642 105472
rect 915 104520 78722 105192
rect 915 104240 78642 104520
rect 915 103568 78722 104240
rect 915 103288 78642 103568
rect 915 102752 78722 103288
rect 915 102472 78642 102752
rect 915 101800 78722 102472
rect 915 101520 78642 101800
rect 915 100848 78722 101520
rect 915 100568 78642 100848
rect 915 99896 78722 100568
rect 915 99616 78642 99896
rect 915 98944 78722 99616
rect 915 98664 78642 98944
rect 915 97992 78722 98664
rect 915 97712 78642 97992
rect 915 97040 78722 97712
rect 915 96760 78642 97040
rect 915 96088 78722 96760
rect 915 95808 78642 96088
rect 915 95136 78722 95808
rect 915 94856 78642 95136
rect 915 94320 78722 94856
rect 915 94040 78642 94320
rect 915 93368 78722 94040
rect 915 93088 78642 93368
rect 915 92416 78722 93088
rect 915 92136 78642 92416
rect 915 91464 78722 92136
rect 915 91184 78642 91464
rect 915 90512 78722 91184
rect 915 90232 78642 90512
rect 915 89560 78722 90232
rect 915 89280 78642 89560
rect 915 88608 78722 89280
rect 915 88328 78642 88608
rect 915 87656 78722 88328
rect 915 87376 78642 87656
rect 915 86704 78722 87376
rect 915 86424 78642 86704
rect 915 85888 78722 86424
rect 915 85608 78642 85888
rect 915 84936 78722 85608
rect 915 84656 78642 84936
rect 915 83984 78722 84656
rect 915 83704 78642 83984
rect 915 83032 78722 83704
rect 915 82752 78642 83032
rect 915 82080 78722 82752
rect 915 81800 78642 82080
rect 915 81128 78722 81800
rect 915 80848 78642 81128
rect 915 80176 78722 80848
rect 915 79896 78642 80176
rect 915 79224 78722 79896
rect 915 78944 78642 79224
rect 915 78272 78722 78944
rect 915 77992 78642 78272
rect 915 77456 78722 77992
rect 915 77176 78642 77456
rect 915 76504 78722 77176
rect 915 76224 78642 76504
rect 915 75552 78722 76224
rect 915 75272 78642 75552
rect 915 74600 78722 75272
rect 915 74320 78642 74600
rect 915 73648 78722 74320
rect 915 73368 78642 73648
rect 915 72696 78722 73368
rect 915 72416 78642 72696
rect 915 71744 78722 72416
rect 915 71464 78642 71744
rect 915 70792 78722 71464
rect 915 70512 78642 70792
rect 915 69840 78722 70512
rect 915 69560 78642 69840
rect 915 69024 78722 69560
rect 915 68744 78642 69024
rect 915 68072 78722 68744
rect 915 67792 78642 68072
rect 915 67120 78722 67792
rect 915 66840 78642 67120
rect 915 66168 78722 66840
rect 915 65888 78642 66168
rect 915 65216 78722 65888
rect 915 64936 78642 65216
rect 915 64264 78722 64936
rect 915 63984 78642 64264
rect 915 63312 78722 63984
rect 915 63032 78642 63312
rect 915 62360 78722 63032
rect 915 62080 78642 62360
rect 915 61408 78722 62080
rect 915 61128 78642 61408
rect 915 60592 78722 61128
rect 915 60312 78642 60592
rect 915 59640 78722 60312
rect 915 59360 78642 59640
rect 915 58688 78722 59360
rect 915 58408 78642 58688
rect 915 57736 78722 58408
rect 915 57456 78642 57736
rect 915 56784 78722 57456
rect 915 56504 78642 56784
rect 915 55832 78722 56504
rect 915 55552 78642 55832
rect 915 54880 78722 55552
rect 915 54600 78642 54880
rect 915 53928 78722 54600
rect 915 53648 78642 53928
rect 915 52976 78722 53648
rect 915 52696 78642 52976
rect 915 52024 78722 52696
rect 915 51744 78642 52024
rect 915 51208 78722 51744
rect 915 50928 78642 51208
rect 915 50256 78722 50928
rect 915 49976 78642 50256
rect 915 49304 78722 49976
rect 915 49024 78642 49304
rect 915 48352 78722 49024
rect 915 48072 78642 48352
rect 915 47400 78722 48072
rect 915 47120 78642 47400
rect 915 46448 78722 47120
rect 915 46168 78642 46448
rect 915 45496 78722 46168
rect 915 45216 78642 45496
rect 915 44544 78722 45216
rect 915 44264 78642 44544
rect 915 43592 78722 44264
rect 915 43312 78642 43592
rect 915 42776 78722 43312
rect 915 42496 78642 42776
rect 915 41824 78722 42496
rect 915 41544 78642 41824
rect 915 40872 78722 41544
rect 915 40592 78642 40872
rect 915 39920 78722 40592
rect 915 39640 78642 39920
rect 915 38968 78722 39640
rect 915 38688 78642 38968
rect 915 38016 78722 38688
rect 915 37736 78642 38016
rect 915 37064 78722 37736
rect 915 36784 78642 37064
rect 915 36112 78722 36784
rect 915 35832 78642 36112
rect 915 35160 78722 35832
rect 915 34880 78642 35160
rect 915 34344 78722 34880
rect 915 34064 78642 34344
rect 915 33392 78722 34064
rect 915 33112 78642 33392
rect 915 32440 78722 33112
rect 915 32160 78642 32440
rect 915 31488 78722 32160
rect 915 31208 78642 31488
rect 915 30536 78722 31208
rect 915 30256 78642 30536
rect 915 29584 78722 30256
rect 915 29304 78642 29584
rect 915 28632 78722 29304
rect 915 28352 78642 28632
rect 915 27680 78722 28352
rect 915 27400 78642 27680
rect 915 26728 78722 27400
rect 915 26448 78642 26728
rect 915 25912 78722 26448
rect 915 25632 78642 25912
rect 915 24960 78722 25632
rect 915 24680 78642 24960
rect 915 24008 78722 24680
rect 915 23728 78642 24008
rect 915 23056 78722 23728
rect 915 22776 78642 23056
rect 915 22104 78722 22776
rect 915 21824 78642 22104
rect 915 21152 78722 21824
rect 915 20872 78642 21152
rect 915 20200 78722 20872
rect 915 19920 78642 20200
rect 915 19248 78722 19920
rect 915 18968 78642 19248
rect 915 18296 78722 18968
rect 915 18016 78642 18296
rect 915 17480 78722 18016
rect 915 17200 78642 17480
rect 915 16528 78722 17200
rect 915 16248 78642 16528
rect 915 15576 78722 16248
rect 915 15296 78642 15576
rect 915 14624 78722 15296
rect 915 14344 78642 14624
rect 915 13672 78722 14344
rect 915 13392 78642 13672
rect 915 12720 78722 13392
rect 915 12440 78642 12720
rect 915 11768 78722 12440
rect 915 11488 78642 11768
rect 915 10816 78722 11488
rect 915 10536 78642 10816
rect 915 9864 78722 10536
rect 915 9584 78642 9864
rect 915 9048 78722 9584
rect 915 8768 78642 9048
rect 915 8096 78722 8768
rect 915 7816 78642 8096
rect 915 7144 78722 7816
rect 915 6864 78642 7144
rect 915 6192 78722 6864
rect 915 5912 78642 6192
rect 915 5240 78722 5912
rect 915 4960 78642 5240
rect 915 4288 78722 4960
rect 915 4008 78642 4288
rect 915 3336 78722 4008
rect 915 3056 78642 3336
rect 915 2384 78722 3056
rect 915 2104 78642 2384
rect 915 1432 78722 2104
rect 915 1152 78642 1432
rect 915 616 78722 1152
rect 915 443 78642 616
<< metal4 >>
rect 3730 2128 4050 117552
rect 19090 2128 19410 117552
rect 34450 2128 34770 117552
rect 49810 2128 50130 117552
rect 65170 2128 65490 117552
<< obsm4 >>
rect 9149 3435 19010 115157
rect 19490 3435 34370 115157
rect 34850 3435 49730 115157
rect 50210 3435 65090 115157
rect 65570 3435 76927 115157
<< labels >>
rlabel metal2 s 0 119200 56 120000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 9936 119200 9992 120000 6 A[10]
port 2 nsew signal input
rlabel metal2 s 10948 119200 11004 120000 6 A[11]
port 3 nsew signal input
rlabel metal2 s 11960 119200 12016 120000 6 A[12]
port 4 nsew signal input
rlabel metal2 s 12972 119200 13028 120000 6 A[13]
port 5 nsew signal input
rlabel metal2 s 13984 119200 14040 120000 6 A[14]
port 6 nsew signal input
rlabel metal2 s 14996 119200 15052 120000 6 A[15]
port 7 nsew signal input
rlabel metal2 s 16008 119200 16064 120000 6 A[16]
port 8 nsew signal input
rlabel metal2 s 16928 119200 16984 120000 6 A[17]
port 9 nsew signal input
rlabel metal2 s 17940 119200 17996 120000 6 A[18]
port 10 nsew signal input
rlabel metal2 s 18952 119200 19008 120000 6 A[19]
port 11 nsew signal input
rlabel metal2 s 920 119200 976 120000 6 A[1]
port 12 nsew signal input
rlabel metal2 s 19964 119200 20020 120000 6 A[20]
port 13 nsew signal input
rlabel metal2 s 20976 119200 21032 120000 6 A[21]
port 14 nsew signal input
rlabel metal2 s 21988 119200 22044 120000 6 A[22]
port 15 nsew signal input
rlabel metal2 s 23000 119200 23056 120000 6 A[23]
port 16 nsew signal input
rlabel metal2 s 1932 119200 1988 120000 6 A[2]
port 17 nsew signal input
rlabel metal2 s 2944 119200 3000 120000 6 A[3]
port 18 nsew signal input
rlabel metal2 s 3956 119200 4012 120000 6 A[4]
port 19 nsew signal input
rlabel metal2 s 4968 119200 5024 120000 6 A[5]
port 20 nsew signal input
rlabel metal2 s 5980 119200 6036 120000 6 A[6]
port 21 nsew signal input
rlabel metal2 s 6992 119200 7048 120000 6 A[7]
port 22 nsew signal input
rlabel metal2 s 8004 119200 8060 120000 6 A[8]
port 23 nsew signal input
rlabel metal2 s 8924 119200 8980 120000 6 A[9]
port 24 nsew signal input
rlabel metal2 s 24012 119200 24068 120000 6 A_h[0]
port 25 nsew signal input
rlabel metal2 s 33948 119200 34004 120000 6 A_h[10]
port 26 nsew signal input
rlabel metal2 s 34960 119200 35016 120000 6 A_h[11]
port 27 nsew signal input
rlabel metal2 s 35972 119200 36028 120000 6 A_h[12]
port 28 nsew signal input
rlabel metal2 s 36984 119200 37040 120000 6 A_h[13]
port 29 nsew signal input
rlabel metal2 s 37996 119200 38052 120000 6 A_h[14]
port 30 nsew signal input
rlabel metal2 s 39008 119200 39064 120000 6 A_h[15]
port 31 nsew signal input
rlabel metal2 s 40020 119200 40076 120000 6 A_h[16]
port 32 nsew signal input
rlabel metal2 s 40940 119200 40996 120000 6 A_h[17]
port 33 nsew signal input
rlabel metal2 s 41952 119200 42008 120000 6 A_h[18]
port 34 nsew signal input
rlabel metal2 s 42964 119200 43020 120000 6 A_h[19]
port 35 nsew signal input
rlabel metal2 s 24932 119200 24988 120000 6 A_h[1]
port 36 nsew signal input
rlabel metal2 s 43976 119200 44032 120000 6 A_h[20]
port 37 nsew signal input
rlabel metal2 s 44988 119200 45044 120000 6 A_h[21]
port 38 nsew signal input
rlabel metal2 s 46000 119200 46056 120000 6 A_h[22]
port 39 nsew signal input
rlabel metal2 s 47012 119200 47068 120000 6 A_h[23]
port 40 nsew signal input
rlabel metal2 s 25944 119200 26000 120000 6 A_h[2]
port 41 nsew signal input
rlabel metal2 s 26956 119200 27012 120000 6 A_h[3]
port 42 nsew signal input
rlabel metal2 s 27968 119200 28024 120000 6 A_h[4]
port 43 nsew signal input
rlabel metal2 s 28980 119200 29036 120000 6 A_h[5]
port 44 nsew signal input
rlabel metal2 s 29992 119200 30048 120000 6 A_h[6]
port 45 nsew signal input
rlabel metal2 s 31004 119200 31060 120000 6 A_h[7]
port 46 nsew signal input
rlabel metal2 s 32016 119200 32072 120000 6 A_h[8]
port 47 nsew signal input
rlabel metal2 s 32936 119200 32992 120000 6 A_h[9]
port 48 nsew signal input
rlabel metal2 s 48024 119200 48080 120000 6 Do[0]
port 49 nsew signal output
rlabel metal2 s 57960 119200 58016 120000 6 Do[10]
port 50 nsew signal output
rlabel metal2 s 58972 119200 59028 120000 6 Do[11]
port 51 nsew signal output
rlabel metal2 s 59984 119200 60040 120000 6 Do[12]
port 52 nsew signal output
rlabel metal2 s 60996 119200 61052 120000 6 Do[13]
port 53 nsew signal output
rlabel metal2 s 62008 119200 62064 120000 6 Do[14]
port 54 nsew signal output
rlabel metal2 s 63020 119200 63076 120000 6 Do[15]
port 55 nsew signal output
rlabel metal2 s 64032 119200 64088 120000 6 Do[16]
port 56 nsew signal output
rlabel metal2 s 64952 119200 65008 120000 6 Do[17]
port 57 nsew signal output
rlabel metal2 s 65964 119200 66020 120000 6 Do[18]
port 58 nsew signal output
rlabel metal2 s 66976 119200 67032 120000 6 Do[19]
port 59 nsew signal output
rlabel metal2 s 48944 119200 49000 120000 6 Do[1]
port 60 nsew signal output
rlabel metal2 s 67988 119200 68044 120000 6 Do[20]
port 61 nsew signal output
rlabel metal2 s 69000 119200 69056 120000 6 Do[21]
port 62 nsew signal output
rlabel metal2 s 70012 119200 70068 120000 6 Do[22]
port 63 nsew signal output
rlabel metal2 s 71024 119200 71080 120000 6 Do[23]
port 64 nsew signal output
rlabel metal2 s 72036 119200 72092 120000 6 Do[24]
port 65 nsew signal output
rlabel metal2 s 72956 119200 73012 120000 6 Do[25]
port 66 nsew signal output
rlabel metal2 s 73968 119200 74024 120000 6 Do[26]
port 67 nsew signal output
rlabel metal2 s 74980 119200 75036 120000 6 Do[27]
port 68 nsew signal output
rlabel metal2 s 75992 119200 76048 120000 6 Do[28]
port 69 nsew signal output
rlabel metal2 s 77004 119200 77060 120000 6 Do[29]
port 70 nsew signal output
rlabel metal2 s 49956 119200 50012 120000 6 Do[2]
port 71 nsew signal output
rlabel metal2 s 78016 119200 78072 120000 6 Do[30]
port 72 nsew signal output
rlabel metal2 s 79028 119200 79084 120000 6 Do[31]
port 73 nsew signal output
rlabel metal2 s 50968 119200 51024 120000 6 Do[3]
port 74 nsew signal output
rlabel metal2 s 51980 119200 52036 120000 6 Do[4]
port 75 nsew signal output
rlabel metal2 s 52992 119200 53048 120000 6 Do[5]
port 76 nsew signal output
rlabel metal2 s 54004 119200 54060 120000 6 Do[6]
port 77 nsew signal output
rlabel metal2 s 55016 119200 55072 120000 6 Do[7]
port 78 nsew signal output
rlabel metal2 s 56028 119200 56084 120000 6 Do[8]
port 79 nsew signal output
rlabel metal2 s 56948 119200 57004 120000 6 Do[9]
port 80 nsew signal output
rlabel metal2 s 9476 0 9532 800 6 clk
port 81 nsew signal input
rlabel metal2 s 69460 0 69516 800 6 hit
port 82 nsew signal output
rlabel metal3 s 78722 416 79522 536 6 line[0]
port 83 nsew signal input
rlabel metal3 s 78722 94120 79522 94240 6 line[100]
port 84 nsew signal input
rlabel metal3 s 78722 94936 79522 95056 6 line[101]
port 85 nsew signal input
rlabel metal3 s 78722 95888 79522 96008 6 line[102]
port 86 nsew signal input
rlabel metal3 s 78722 96840 79522 96960 6 line[103]
port 87 nsew signal input
rlabel metal3 s 78722 97792 79522 97912 6 line[104]
port 88 nsew signal input
rlabel metal3 s 78722 98744 79522 98864 6 line[105]
port 89 nsew signal input
rlabel metal3 s 78722 99696 79522 99816 6 line[106]
port 90 nsew signal input
rlabel metal3 s 78722 100648 79522 100768 6 line[107]
port 91 nsew signal input
rlabel metal3 s 78722 101600 79522 101720 6 line[108]
port 92 nsew signal input
rlabel metal3 s 78722 102552 79522 102672 6 line[109]
port 93 nsew signal input
rlabel metal3 s 78722 9664 79522 9784 6 line[10]
port 94 nsew signal input
rlabel metal3 s 78722 103368 79522 103488 6 line[110]
port 95 nsew signal input
rlabel metal3 s 78722 104320 79522 104440 6 line[111]
port 96 nsew signal input
rlabel metal3 s 78722 105272 79522 105392 6 line[112]
port 97 nsew signal input
rlabel metal3 s 78722 106224 79522 106344 6 line[113]
port 98 nsew signal input
rlabel metal3 s 78722 107176 79522 107296 6 line[114]
port 99 nsew signal input
rlabel metal3 s 78722 108128 79522 108248 6 line[115]
port 100 nsew signal input
rlabel metal3 s 78722 109080 79522 109200 6 line[116]
port 101 nsew signal input
rlabel metal3 s 78722 110032 79522 110152 6 line[117]
port 102 nsew signal input
rlabel metal3 s 78722 110984 79522 111104 6 line[118]
port 103 nsew signal input
rlabel metal3 s 78722 111800 79522 111920 6 line[119]
port 104 nsew signal input
rlabel metal3 s 78722 10616 79522 10736 6 line[11]
port 105 nsew signal input
rlabel metal3 s 78722 112752 79522 112872 6 line[120]
port 106 nsew signal input
rlabel metal3 s 78722 113704 79522 113824 6 line[121]
port 107 nsew signal input
rlabel metal3 s 78722 114656 79522 114776 6 line[122]
port 108 nsew signal input
rlabel metal3 s 78722 115608 79522 115728 6 line[123]
port 109 nsew signal input
rlabel metal3 s 78722 116560 79522 116680 6 line[124]
port 110 nsew signal input
rlabel metal3 s 78722 117512 79522 117632 6 line[125]
port 111 nsew signal input
rlabel metal3 s 78722 118464 79522 118584 6 line[126]
port 112 nsew signal input
rlabel metal3 s 78722 119416 79522 119536 6 line[127]
port 113 nsew signal input
rlabel metal3 s 78722 11568 79522 11688 6 line[12]
port 114 nsew signal input
rlabel metal3 s 78722 12520 79522 12640 6 line[13]
port 115 nsew signal input
rlabel metal3 s 78722 13472 79522 13592 6 line[14]
port 116 nsew signal input
rlabel metal3 s 78722 14424 79522 14544 6 line[15]
port 117 nsew signal input
rlabel metal3 s 78722 15376 79522 15496 6 line[16]
port 118 nsew signal input
rlabel metal3 s 78722 16328 79522 16448 6 line[17]
port 119 nsew signal input
rlabel metal3 s 78722 17280 79522 17400 6 line[18]
port 120 nsew signal input
rlabel metal3 s 78722 18096 79522 18216 6 line[19]
port 121 nsew signal input
rlabel metal3 s 78722 1232 79522 1352 6 line[1]
port 122 nsew signal input
rlabel metal3 s 78722 19048 79522 19168 6 line[20]
port 123 nsew signal input
rlabel metal3 s 78722 20000 79522 20120 6 line[21]
port 124 nsew signal input
rlabel metal3 s 78722 20952 79522 21072 6 line[22]
port 125 nsew signal input
rlabel metal3 s 78722 21904 79522 22024 6 line[23]
port 126 nsew signal input
rlabel metal3 s 78722 22856 79522 22976 6 line[24]
port 127 nsew signal input
rlabel metal3 s 78722 23808 79522 23928 6 line[25]
port 128 nsew signal input
rlabel metal3 s 78722 24760 79522 24880 6 line[26]
port 129 nsew signal input
rlabel metal3 s 78722 25712 79522 25832 6 line[27]
port 130 nsew signal input
rlabel metal3 s 78722 26528 79522 26648 6 line[28]
port 131 nsew signal input
rlabel metal3 s 78722 27480 79522 27600 6 line[29]
port 132 nsew signal input
rlabel metal3 s 78722 2184 79522 2304 6 line[2]
port 133 nsew signal input
rlabel metal3 s 78722 28432 79522 28552 6 line[30]
port 134 nsew signal input
rlabel metal3 s 78722 29384 79522 29504 6 line[31]
port 135 nsew signal input
rlabel metal3 s 78722 30336 79522 30456 6 line[32]
port 136 nsew signal input
rlabel metal3 s 78722 31288 79522 31408 6 line[33]
port 137 nsew signal input
rlabel metal3 s 78722 32240 79522 32360 6 line[34]
port 138 nsew signal input
rlabel metal3 s 78722 33192 79522 33312 6 line[35]
port 139 nsew signal input
rlabel metal3 s 78722 34144 79522 34264 6 line[36]
port 140 nsew signal input
rlabel metal3 s 78722 34960 79522 35080 6 line[37]
port 141 nsew signal input
rlabel metal3 s 78722 35912 79522 36032 6 line[38]
port 142 nsew signal input
rlabel metal3 s 78722 36864 79522 36984 6 line[39]
port 143 nsew signal input
rlabel metal3 s 78722 3136 79522 3256 6 line[3]
port 144 nsew signal input
rlabel metal3 s 78722 37816 79522 37936 6 line[40]
port 145 nsew signal input
rlabel metal3 s 78722 38768 79522 38888 6 line[41]
port 146 nsew signal input
rlabel metal3 s 78722 39720 79522 39840 6 line[42]
port 147 nsew signal input
rlabel metal3 s 78722 40672 79522 40792 6 line[43]
port 148 nsew signal input
rlabel metal3 s 78722 41624 79522 41744 6 line[44]
port 149 nsew signal input
rlabel metal3 s 78722 42576 79522 42696 6 line[45]
port 150 nsew signal input
rlabel metal3 s 78722 43392 79522 43512 6 line[46]
port 151 nsew signal input
rlabel metal3 s 78722 44344 79522 44464 6 line[47]
port 152 nsew signal input
rlabel metal3 s 78722 45296 79522 45416 6 line[48]
port 153 nsew signal input
rlabel metal3 s 78722 46248 79522 46368 6 line[49]
port 154 nsew signal input
rlabel metal3 s 78722 4088 79522 4208 6 line[4]
port 155 nsew signal input
rlabel metal3 s 78722 47200 79522 47320 6 line[50]
port 156 nsew signal input
rlabel metal3 s 78722 48152 79522 48272 6 line[51]
port 157 nsew signal input
rlabel metal3 s 78722 49104 79522 49224 6 line[52]
port 158 nsew signal input
rlabel metal3 s 78722 50056 79522 50176 6 line[53]
port 159 nsew signal input
rlabel metal3 s 78722 51008 79522 51128 6 line[54]
port 160 nsew signal input
rlabel metal3 s 78722 51824 79522 51944 6 line[55]
port 161 nsew signal input
rlabel metal3 s 78722 52776 79522 52896 6 line[56]
port 162 nsew signal input
rlabel metal3 s 78722 53728 79522 53848 6 line[57]
port 163 nsew signal input
rlabel metal3 s 78722 54680 79522 54800 6 line[58]
port 164 nsew signal input
rlabel metal3 s 78722 55632 79522 55752 6 line[59]
port 165 nsew signal input
rlabel metal3 s 78722 5040 79522 5160 6 line[5]
port 166 nsew signal input
rlabel metal3 s 78722 56584 79522 56704 6 line[60]
port 167 nsew signal input
rlabel metal3 s 78722 57536 79522 57656 6 line[61]
port 168 nsew signal input
rlabel metal3 s 78722 58488 79522 58608 6 line[62]
port 169 nsew signal input
rlabel metal3 s 78722 59440 79522 59560 6 line[63]
port 170 nsew signal input
rlabel metal3 s 78722 60392 79522 60512 6 line[64]
port 171 nsew signal input
rlabel metal3 s 78722 61208 79522 61328 6 line[65]
port 172 nsew signal input
rlabel metal3 s 78722 62160 79522 62280 6 line[66]
port 173 nsew signal input
rlabel metal3 s 78722 63112 79522 63232 6 line[67]
port 174 nsew signal input
rlabel metal3 s 78722 64064 79522 64184 6 line[68]
port 175 nsew signal input
rlabel metal3 s 78722 65016 79522 65136 6 line[69]
port 176 nsew signal input
rlabel metal3 s 78722 5992 79522 6112 6 line[6]
port 177 nsew signal input
rlabel metal3 s 78722 65968 79522 66088 6 line[70]
port 178 nsew signal input
rlabel metal3 s 78722 66920 79522 67040 6 line[71]
port 179 nsew signal input
rlabel metal3 s 78722 67872 79522 67992 6 line[72]
port 180 nsew signal input
rlabel metal3 s 78722 68824 79522 68944 6 line[73]
port 181 nsew signal input
rlabel metal3 s 78722 69640 79522 69760 6 line[74]
port 182 nsew signal input
rlabel metal3 s 78722 70592 79522 70712 6 line[75]
port 183 nsew signal input
rlabel metal3 s 78722 71544 79522 71664 6 line[76]
port 184 nsew signal input
rlabel metal3 s 78722 72496 79522 72616 6 line[77]
port 185 nsew signal input
rlabel metal3 s 78722 73448 79522 73568 6 line[78]
port 186 nsew signal input
rlabel metal3 s 78722 74400 79522 74520 6 line[79]
port 187 nsew signal input
rlabel metal3 s 78722 6944 79522 7064 6 line[7]
port 188 nsew signal input
rlabel metal3 s 78722 75352 79522 75472 6 line[80]
port 189 nsew signal input
rlabel metal3 s 78722 76304 79522 76424 6 line[81]
port 190 nsew signal input
rlabel metal3 s 78722 77256 79522 77376 6 line[82]
port 191 nsew signal input
rlabel metal3 s 78722 78072 79522 78192 6 line[83]
port 192 nsew signal input
rlabel metal3 s 78722 79024 79522 79144 6 line[84]
port 193 nsew signal input
rlabel metal3 s 78722 79976 79522 80096 6 line[85]
port 194 nsew signal input
rlabel metal3 s 78722 80928 79522 81048 6 line[86]
port 195 nsew signal input
rlabel metal3 s 78722 81880 79522 82000 6 line[87]
port 196 nsew signal input
rlabel metal3 s 78722 82832 79522 82952 6 line[88]
port 197 nsew signal input
rlabel metal3 s 78722 83784 79522 83904 6 line[89]
port 198 nsew signal input
rlabel metal3 s 78722 7896 79522 8016 6 line[8]
port 199 nsew signal input
rlabel metal3 s 78722 84736 79522 84856 6 line[90]
port 200 nsew signal input
rlabel metal3 s 78722 85688 79522 85808 6 line[91]
port 201 nsew signal input
rlabel metal3 s 78722 86504 79522 86624 6 line[92]
port 202 nsew signal input
rlabel metal3 s 78722 87456 79522 87576 6 line[93]
port 203 nsew signal input
rlabel metal3 s 78722 88408 79522 88528 6 line[94]
port 204 nsew signal input
rlabel metal3 s 78722 89360 79522 89480 6 line[95]
port 205 nsew signal input
rlabel metal3 s 78722 90312 79522 90432 6 line[96]
port 206 nsew signal input
rlabel metal3 s 78722 91264 79522 91384 6 line[97]
port 207 nsew signal input
rlabel metal3 s 78722 92216 79522 92336 6 line[98]
port 208 nsew signal input
rlabel metal3 s 78722 93168 79522 93288 6 line[99]
port 209 nsew signal input
rlabel metal3 s 78722 8848 79522 8968 6 line[9]
port 210 nsew signal input
rlabel metal2 s 29440 0 29496 800 6 rst_n
port 211 nsew signal input
rlabel metal2 s 49496 0 49552 800 6 wr
port 212 nsew signal input
rlabel metal4 s 65170 2128 65490 117552 6 VPWR
port 213 nsew power bidirectional
rlabel metal4 s 34450 2128 34770 117552 6 VPWR
port 214 nsew power bidirectional
rlabel metal4 s 3730 2128 4050 117552 6 VPWR
port 215 nsew power bidirectional
rlabel metal4 s 49810 2128 50130 117552 6 VGND
port 216 nsew ground bidirectional
rlabel metal4 s 19090 2128 19410 117552 6 VGND
port 217 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 79522 120000
string LEFview TRUE
<< end >>
