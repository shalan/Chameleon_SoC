magic
tech sky130A
magscale 1 2
timestamp 1608830673
<< obsli1 >>
rect 38 31 217802 275329
<< obsm1 >>
rect 38 0 217802 275440
<< metal2 >>
rect 332 277072 388 277872
rect 3092 277072 3148 277872
rect 5944 277072 6000 277872
rect 8704 277072 8760 277872
rect 11556 277072 11612 277872
rect 14408 277072 14464 277872
rect 17168 277072 17224 277872
rect 20020 277072 20076 277872
rect 22872 277072 22928 277872
rect 25632 277072 25688 277872
rect 28484 277072 28540 277872
rect 31336 277072 31392 277872
rect 34096 277072 34152 277872
rect 36948 277072 37004 277872
rect 39800 277072 39856 277872
rect 42560 277072 42616 277872
rect 45412 277072 45468 277872
rect 48264 277072 48320 277872
rect 51024 277072 51080 277872
rect 53876 277072 53932 277872
rect 56728 277072 56784 277872
rect 59488 277072 59544 277872
rect 62340 277072 62396 277872
rect 65192 277072 65248 277872
rect 67952 277072 68008 277872
rect 70804 277072 70860 277872
rect 73656 277072 73712 277872
rect 76416 277072 76472 277872
rect 79268 277072 79324 277872
rect 82028 277072 82084 277872
rect 84880 277072 84936 277872
rect 87732 277072 87788 277872
rect 90492 277072 90548 277872
rect 93344 277072 93400 277872
rect 96196 277072 96252 277872
rect 98956 277072 99012 277872
rect 101808 277072 101864 277872
rect 104660 277072 104716 277872
rect 107420 277072 107476 277872
rect 110272 277072 110328 277872
rect 113124 277072 113180 277872
rect 115884 277072 115940 277872
rect 118736 277072 118792 277872
rect 121588 277072 121644 277872
rect 124348 277072 124404 277872
rect 127200 277072 127256 277872
rect 130052 277072 130108 277872
rect 132812 277072 132868 277872
rect 135664 277072 135720 277872
rect 138516 277072 138572 277872
rect 141276 277072 141332 277872
rect 144128 277072 144184 277872
rect 146980 277072 147036 277872
rect 149740 277072 149796 277872
rect 152592 277072 152648 277872
rect 155352 277072 155408 277872
rect 158204 277072 158260 277872
rect 161056 277072 161112 277872
rect 163816 277072 163872 277872
rect 166668 277072 166724 277872
rect 169520 277072 169576 277872
rect 172280 277072 172336 277872
rect 175132 277072 175188 277872
rect 177984 277072 178040 277872
rect 180744 277072 180800 277872
rect 183596 277072 183652 277872
rect 186448 277072 186504 277872
rect 189208 277072 189264 277872
rect 192060 277072 192116 277872
rect 194912 277072 194968 277872
rect 197672 277072 197728 277872
rect 200524 277072 200580 277872
rect 203376 277072 203432 277872
rect 206136 277072 206192 277872
rect 208988 277072 209044 277872
rect 211840 277072 211896 277872
rect 214600 277072 214656 277872
rect 217452 277072 217508 277872
<< obsm2 >>
rect 444 277016 3036 277072
rect 3204 277016 5888 277072
rect 6056 277016 8648 277072
rect 8816 277016 11500 277072
rect 11668 277016 14352 277072
rect 14520 277016 17112 277072
rect 17280 277016 19964 277072
rect 20132 277016 22816 277072
rect 22984 277016 25576 277072
rect 25744 277016 28428 277072
rect 28596 277016 31280 277072
rect 31448 277016 34040 277072
rect 34208 277016 36892 277072
rect 37060 277016 39744 277072
rect 39912 277016 42504 277072
rect 42672 277016 45356 277072
rect 45524 277016 48208 277072
rect 48376 277016 50968 277072
rect 51136 277016 53820 277072
rect 53988 277016 56672 277072
rect 56840 277016 59432 277072
rect 59600 277016 62284 277072
rect 62452 277016 65136 277072
rect 65304 277016 67896 277072
rect 68064 277016 70748 277072
rect 70916 277016 73600 277072
rect 73768 277016 76360 277072
rect 76528 277016 79212 277072
rect 79380 277016 81972 277072
rect 82140 277016 84824 277072
rect 84992 277016 87676 277072
rect 87844 277016 90436 277072
rect 90604 277016 93288 277072
rect 93456 277016 96140 277072
rect 96308 277016 98900 277072
rect 99068 277016 101752 277072
rect 101920 277016 104604 277072
rect 104772 277016 107364 277072
rect 107532 277016 110216 277072
rect 110384 277016 113068 277072
rect 113236 277016 115828 277072
rect 115996 277016 118680 277072
rect 118848 277016 121532 277072
rect 121700 277016 124292 277072
rect 124460 277016 127144 277072
rect 127312 277016 129996 277072
rect 130164 277016 132756 277072
rect 132924 277016 135608 277072
rect 135776 277016 138460 277072
rect 138628 277016 141220 277072
rect 141388 277016 144072 277072
rect 144240 277016 146924 277072
rect 147092 277016 149684 277072
rect 149852 277016 152536 277072
rect 152704 277016 155296 277072
rect 155464 277016 158148 277072
rect 158316 277016 161000 277072
rect 161168 277016 163760 277072
rect 163928 277016 166612 277072
rect 166780 277016 169464 277072
rect 169632 277016 172224 277072
rect 172392 277016 175076 277072
rect 175244 277016 177928 277072
rect 178096 277016 180688 277072
rect 180856 277016 183540 277072
rect 183708 277016 186392 277072
rect 186560 277016 189152 277072
rect 189320 277016 192004 277072
rect 192172 277016 194856 277072
rect 195024 277016 197616 277072
rect 197784 277016 200468 277072
rect 200636 277016 203320 277072
rect 203488 277016 206080 277072
rect 206248 277016 208932 277072
rect 209100 277016 211784 277072
rect 211952 277016 214544 277072
rect 214712 277016 217396 277072
rect 334 0 217506 277016
<< obsm3 >>
rect 879 15 203142 275345
<< metal4 >>
rect 3142 0 3462 275360
rect 18502 0 18822 275360
rect 33862 0 34182 275360
rect 49222 0 49542 275360
rect 64582 0 64902 275360
rect 79942 0 80262 275360
rect 95302 0 95622 275360
rect 110662 0 110982 275360
rect 126022 0 126342 275360
rect 141382 0 141702 275360
rect 156742 0 157062 275360
rect 172102 0 172422 275360
rect 187462 0 187782 275360
rect 202822 0 203142 275360
<< obsm4 >>
rect 27881 150635 33782 274869
rect 34262 150635 49142 274869
rect 49622 150635 64502 274869
rect 64982 150635 79862 274869
rect 80342 150635 95222 274869
rect 95702 150635 110582 274869
rect 111062 150635 125942 274869
rect 126422 150635 141302 274869
rect 141782 150635 156662 274869
rect 157142 150635 169259 274869
<< labels >>
rlabel metal2 s 90492 277072 90548 277872 6 A[0]
port 1 nsew signal input
rlabel metal2 s 93344 277072 93400 277872 6 A[1]
port 2 nsew signal input
rlabel metal2 s 96196 277072 96252 277872 6 A[2]
port 3 nsew signal input
rlabel metal2 s 98956 277072 99012 277872 6 A[3]
port 4 nsew signal input
rlabel metal2 s 101808 277072 101864 277872 6 A[4]
port 5 nsew signal input
rlabel metal2 s 104660 277072 104716 277872 6 A[5]
port 6 nsew signal input
rlabel metal2 s 107420 277072 107476 277872 6 A[6]
port 7 nsew signal input
rlabel metal2 s 110272 277072 110328 277872 6 A[7]
port 8 nsew signal input
rlabel metal2 s 113124 277072 113180 277872 6 CLK
port 9 nsew signal input
rlabel metal2 s 130052 277072 130108 277872 6 Di[0]
port 10 nsew signal input
rlabel metal2 s 158204 277072 158260 277872 6 Di[10]
port 11 nsew signal input
rlabel metal2 s 161056 277072 161112 277872 6 Di[11]
port 12 nsew signal input
rlabel metal2 s 163816 277072 163872 277872 6 Di[12]
port 13 nsew signal input
rlabel metal2 s 166668 277072 166724 277872 6 Di[13]
port 14 nsew signal input
rlabel metal2 s 169520 277072 169576 277872 6 Di[14]
port 15 nsew signal input
rlabel metal2 s 172280 277072 172336 277872 6 Di[15]
port 16 nsew signal input
rlabel metal2 s 175132 277072 175188 277872 6 Di[16]
port 17 nsew signal input
rlabel metal2 s 177984 277072 178040 277872 6 Di[17]
port 18 nsew signal input
rlabel metal2 s 180744 277072 180800 277872 6 Di[18]
port 19 nsew signal input
rlabel metal2 s 183596 277072 183652 277872 6 Di[19]
port 20 nsew signal input
rlabel metal2 s 132812 277072 132868 277872 6 Di[1]
port 21 nsew signal input
rlabel metal2 s 186448 277072 186504 277872 6 Di[20]
port 22 nsew signal input
rlabel metal2 s 189208 277072 189264 277872 6 Di[21]
port 23 nsew signal input
rlabel metal2 s 192060 277072 192116 277872 6 Di[22]
port 24 nsew signal input
rlabel metal2 s 194912 277072 194968 277872 6 Di[23]
port 25 nsew signal input
rlabel metal2 s 197672 277072 197728 277872 6 Di[24]
port 26 nsew signal input
rlabel metal2 s 200524 277072 200580 277872 6 Di[25]
port 27 nsew signal input
rlabel metal2 s 203376 277072 203432 277872 6 Di[26]
port 28 nsew signal input
rlabel metal2 s 206136 277072 206192 277872 6 Di[27]
port 29 nsew signal input
rlabel metal2 s 208988 277072 209044 277872 6 Di[28]
port 30 nsew signal input
rlabel metal2 s 211840 277072 211896 277872 6 Di[29]
port 31 nsew signal input
rlabel metal2 s 135664 277072 135720 277872 6 Di[2]
port 32 nsew signal input
rlabel metal2 s 214600 277072 214656 277872 6 Di[30]
port 33 nsew signal input
rlabel metal2 s 217452 277072 217508 277872 6 Di[31]
port 34 nsew signal input
rlabel metal2 s 138516 277072 138572 277872 6 Di[3]
port 35 nsew signal input
rlabel metal2 s 141276 277072 141332 277872 6 Di[4]
port 36 nsew signal input
rlabel metal2 s 144128 277072 144184 277872 6 Di[5]
port 37 nsew signal input
rlabel metal2 s 146980 277072 147036 277872 6 Di[6]
port 38 nsew signal input
rlabel metal2 s 149740 277072 149796 277872 6 Di[7]
port 39 nsew signal input
rlabel metal2 s 152592 277072 152648 277872 6 Di[8]
port 40 nsew signal input
rlabel metal2 s 155352 277072 155408 277872 6 Di[9]
port 41 nsew signal input
rlabel metal2 s 332 277072 388 277872 6 Do[0]
port 42 nsew signal output
rlabel metal2 s 28484 277072 28540 277872 6 Do[10]
port 43 nsew signal output
rlabel metal2 s 31336 277072 31392 277872 6 Do[11]
port 44 nsew signal output
rlabel metal2 s 34096 277072 34152 277872 6 Do[12]
port 45 nsew signal output
rlabel metal2 s 36948 277072 37004 277872 6 Do[13]
port 46 nsew signal output
rlabel metal2 s 39800 277072 39856 277872 6 Do[14]
port 47 nsew signal output
rlabel metal2 s 42560 277072 42616 277872 6 Do[15]
port 48 nsew signal output
rlabel metal2 s 45412 277072 45468 277872 6 Do[16]
port 49 nsew signal output
rlabel metal2 s 48264 277072 48320 277872 6 Do[17]
port 50 nsew signal output
rlabel metal2 s 51024 277072 51080 277872 6 Do[18]
port 51 nsew signal output
rlabel metal2 s 53876 277072 53932 277872 6 Do[19]
port 52 nsew signal output
rlabel metal2 s 3092 277072 3148 277872 6 Do[1]
port 53 nsew signal output
rlabel metal2 s 56728 277072 56784 277872 6 Do[20]
port 54 nsew signal output
rlabel metal2 s 59488 277072 59544 277872 6 Do[21]
port 55 nsew signal output
rlabel metal2 s 62340 277072 62396 277872 6 Do[22]
port 56 nsew signal output
rlabel metal2 s 65192 277072 65248 277872 6 Do[23]
port 57 nsew signal output
rlabel metal2 s 67952 277072 68008 277872 6 Do[24]
port 58 nsew signal output
rlabel metal2 s 70804 277072 70860 277872 6 Do[25]
port 59 nsew signal output
rlabel metal2 s 73656 277072 73712 277872 6 Do[26]
port 60 nsew signal output
rlabel metal2 s 76416 277072 76472 277872 6 Do[27]
port 61 nsew signal output
rlabel metal2 s 79268 277072 79324 277872 6 Do[28]
port 62 nsew signal output
rlabel metal2 s 82028 277072 82084 277872 6 Do[29]
port 63 nsew signal output
rlabel metal2 s 5944 277072 6000 277872 6 Do[2]
port 64 nsew signal output
rlabel metal2 s 84880 277072 84936 277872 6 Do[30]
port 65 nsew signal output
rlabel metal2 s 87732 277072 87788 277872 6 Do[31]
port 66 nsew signal output
rlabel metal2 s 8704 277072 8760 277872 6 Do[3]
port 67 nsew signal output
rlabel metal2 s 11556 277072 11612 277872 6 Do[4]
port 68 nsew signal output
rlabel metal2 s 14408 277072 14464 277872 6 Do[5]
port 69 nsew signal output
rlabel metal2 s 17168 277072 17224 277872 6 Do[6]
port 70 nsew signal output
rlabel metal2 s 20020 277072 20076 277872 6 Do[7]
port 71 nsew signal output
rlabel metal2 s 22872 277072 22928 277872 6 Do[8]
port 72 nsew signal output
rlabel metal2 s 25632 277072 25688 277872 6 Do[9]
port 73 nsew signal output
rlabel metal2 s 127200 277072 127256 277872 6 EN
port 74 nsew signal input
rlabel metal2 s 115884 277072 115940 277872 6 WE[0]
port 75 nsew signal input
rlabel metal2 s 118736 277072 118792 277872 6 WE[1]
port 76 nsew signal input
rlabel metal2 s 121588 277072 121644 277872 6 WE[2]
port 77 nsew signal input
rlabel metal2 s 124348 277072 124404 277872 6 WE[3]
port 78 nsew signal input
rlabel metal4 s 187462 0 187782 275360 6 VPWR
port 79 nsew power bidirectional
rlabel metal4 s 156742 0 157062 275360 6 VPWR
port 80 nsew power bidirectional
rlabel metal4 s 126022 0 126342 275360 6 VPWR
port 81 nsew power bidirectional
rlabel metal4 s 95302 0 95622 275360 6 VPWR
port 82 nsew power bidirectional
rlabel metal4 s 64582 0 64902 275360 6 VPWR
port 83 nsew power bidirectional
rlabel metal4 s 33862 0 34182 275360 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 3142 0 3462 275360 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 202822 0 203142 275360 6 VGND
port 86 nsew ground bidirectional
rlabel metal4 s 172102 0 172422 275360 6 VGND
port 87 nsew ground bidirectional
rlabel metal4 s 141382 0 141702 275360 6 VGND
port 88 nsew ground bidirectional
rlabel metal4 s 110662 0 110982 275360 6 VGND
port 89 nsew ground bidirectional
rlabel metal4 s 79942 0 80262 275360 6 VGND
port 90 nsew ground bidirectional
rlabel metal4 s 49222 0 49542 275360 6 VGND
port 91 nsew ground bidirectional
rlabel metal4 s 18502 0 18822 275360 6 VGND
port 92 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 217840 277872
string LEFview TRUE
<< end >>
